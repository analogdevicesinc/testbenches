// ***************************************************************************
// ***************************************************************************
// Copyright (C) 2014 - 2025 Analog Devices, Inc. All rights reserved.
//
// In this HDL repository, there are many different and unique modules, consisting
// of various HDL (Verilog or VHDL) components. The individual modules are
// developed independently, and may be accompanied by separate and unique license
// terms.
//
// The user should read each of these license terms, and understand the
// freedoms and responsabilities that he or she has by using this source/core.
//
// This core is distributed in the hope that it will be useful, but WITHOUT ANY
// WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR
// A PARTICULAR PURPOSE.
//
// Redistribution and use of source or resulting binaries, with or without modification
// of this file, are permitted under one of the following two license terms:
//
//   1. The GNU General Public License version 2 as published by the
//      Free Software Foundation, which can be found in the top level directory
//      of this repository (LICENSE_GPL2), and also online at:
//      <https://www.gnu.org/licenses/old-licenses/gpl-2.0.html>
//
// OR
//
//   2. An ADI specific BSD license, which can be found in the top level directory
//      of this repository (LICENSE_ADIBSD), and also on-line at:
//      https://github.com/analogdevicesinc/hdl/blob/main/LICENSE_ADIBSD
//      This will allow to generate bit files and not release the source code,
//      as long as it attaches to an ADI device.
//
// ***************************************************************************
// ***************************************************************************
/* Auto generated Register Map */
/* Feb 07 11:48:47 2025 v0.4.1 */

`timescale 1ns/1ps

`ifndef _ADI_REGMAP_DATA_OFFLOAD_PKG_DEFINITIONS_SVH_
`define _ADI_REGMAP_DATA_OFFLOAD_PKG_DEFINITIONS_SVH_

// Help build VIP Interface parameters name
`define ADI_REGMAP_DATA_OFFLOAD_PKG_PARAM_IMPORT(n)  n``.inst.AUTO_BRINGUP, \
  n``.inst.HAS_BYPASS, \
  n``.inst.ID, \
  n``.inst.MEM_SIZE_LOG2, \
  n``.inst.MEM_TYPE, \
  n``.inst.TX_OR_RXN_PATH

`define ADI_REGMAP_DATA_OFFLOAD_PKG_PARAM_DECL int  AUTO_BRINGUP, \
  HAS_BYPASS, \
  ID, \
  MEM_SIZE_LOG2, \
  MEM_TYPE, \
  TX_OR_RXN_PATH

`define ADI_REGMAP_DATA_OFFLOAD_PKG_PARAM_ORDER  AUTO_BRINGUP, \
  HAS_BYPASS, \
  ID, \
  MEM_SIZE_LOG2, \
  MEM_TYPE, \
  TX_OR_RXN_PATH

`endif
