// ***************************************************************************
// ***************************************************************************
// Copyright (C) 2014 - 2024 Analog Devices, Inc. All rights reserved.
//
// In this HDL repository, there are many different and unique modules, consisting
// of various HDL (Verilog or VHDL) components. The individual modules are
// developed independently, and may be accompanied by separate and unique license
// terms.
//
// The user should read each of these license terms, and understand the
// freedoms and responsabilities that he or she has by using this source/core.
//
// This core is distributed in the hope that it will be useful, but WITHOUT ANY
// WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR
// A PARTICULAR PURPOSE.
//
// Redistribution and use of source or resulting binaries, with or without modification
// of this file, are permitted under one of the following two license terms:
//
//   1. The GNU General Public License version 2 as published by the
//      Free Software Foundation, which can be found in the top level directory
//      of this repository (LICENSE_GPL2), and also online at:
//      <https://www.gnu.org/licenses/old-licenses/gpl-2.0.html>
//
// OR
//
//   2. An ADI specific BSD license, which can be found in the top level directory
//      of this repository (LICENSE_ADIBSD), and also on-line at:
//      https://github.com/analogdevicesinc/hdl/blob/main/LICENSE_ADIBSD
//      This will allow to generate bit files and not release the source code,
//      as long as it attaches to an ADI device.
//
// ***************************************************************************
// ***************************************************************************
/* Auto generated Register Map */
/* Thu Mar 28 13:22:23 2024 */

package adi_regmap_dac_pkg;
  import adi_regmap_pkg::*;


/* DAC Common (axi_ad) */

  const reg_t DAC_COMMON_REG_RSTN = '{ 'h0040, "REG_RSTN" , '{
    "CE_N": '{ 2, 2, RW, 'h0 },
    "MMCM_RSTN": '{ 1, 1, RW, 'h0 },
    "RSTN": '{ 0, 0, RW, 'h0 }}};
  `define SET_DAC_COMMON_REG_RSTN_CE_N(x) SetField(DAC_COMMON_REG_RSTN,"CE_N",x)
  `define GET_DAC_COMMON_REG_RSTN_CE_N(x) GetField(DAC_COMMON_REG_RSTN,"CE_N",x)
  `define DEFAULT_DAC_COMMON_REG_RSTN_CE_N GetResetValue(DAC_COMMON_REG_RSTN,"CE_N")
  `define UPDATE_DAC_COMMON_REG_RSTN_CE_N(x,y) UpdateField(DAC_COMMON_REG_RSTN,"CE_N",x,y)
  `define SET_DAC_COMMON_REG_RSTN_MMCM_RSTN(x) SetField(DAC_COMMON_REG_RSTN,"MMCM_RSTN",x)
  `define GET_DAC_COMMON_REG_RSTN_MMCM_RSTN(x) GetField(DAC_COMMON_REG_RSTN,"MMCM_RSTN",x)
  `define DEFAULT_DAC_COMMON_REG_RSTN_MMCM_RSTN GetResetValue(DAC_COMMON_REG_RSTN,"MMCM_RSTN")
  `define UPDATE_DAC_COMMON_REG_RSTN_MMCM_RSTN(x,y) UpdateField(DAC_COMMON_REG_RSTN,"MMCM_RSTN",x,y)
  `define SET_DAC_COMMON_REG_RSTN_RSTN(x) SetField(DAC_COMMON_REG_RSTN,"RSTN",x)
  `define GET_DAC_COMMON_REG_RSTN_RSTN(x) GetField(DAC_COMMON_REG_RSTN,"RSTN",x)
  `define DEFAULT_DAC_COMMON_REG_RSTN_RSTN GetResetValue(DAC_COMMON_REG_RSTN,"RSTN")
  `define UPDATE_DAC_COMMON_REG_RSTN_RSTN(x,y) UpdateField(DAC_COMMON_REG_RSTN,"RSTN",x,y)

  const reg_t DAC_COMMON_REG_CNTRL_1 = '{ 'h0044, "REG_CNTRL_1" , '{
    "SYNC": '{ 0, 0, RW, 'h0 },
    "EXT_SYNC_ARM": '{ 1, 1, RW, 'h0 },
    "EXT_SYNC_DISARM": '{ 2, 2, RW, 'h0 },
    "MANUAL_SYNC_REQUEST": '{ 8, 8, RW, 'h0 }}};
  `define SET_DAC_COMMON_REG_CNTRL_1_SYNC(x) SetField(DAC_COMMON_REG_CNTRL_1,"SYNC",x)
  `define GET_DAC_COMMON_REG_CNTRL_1_SYNC(x) GetField(DAC_COMMON_REG_CNTRL_1,"SYNC",x)
  `define DEFAULT_DAC_COMMON_REG_CNTRL_1_SYNC GetResetValue(DAC_COMMON_REG_CNTRL_1,"SYNC")
  `define UPDATE_DAC_COMMON_REG_CNTRL_1_SYNC(x,y) UpdateField(DAC_COMMON_REG_CNTRL_1,"SYNC",x,y)
  `define SET_DAC_COMMON_REG_CNTRL_1_EXT_SYNC_ARM(x) SetField(DAC_COMMON_REG_CNTRL_1,"EXT_SYNC_ARM",x)
  `define GET_DAC_COMMON_REG_CNTRL_1_EXT_SYNC_ARM(x) GetField(DAC_COMMON_REG_CNTRL_1,"EXT_SYNC_ARM",x)
  `define DEFAULT_DAC_COMMON_REG_CNTRL_1_EXT_SYNC_ARM GetResetValue(DAC_COMMON_REG_CNTRL_1,"EXT_SYNC_ARM")
  `define UPDATE_DAC_COMMON_REG_CNTRL_1_EXT_SYNC_ARM(x,y) UpdateField(DAC_COMMON_REG_CNTRL_1,"EXT_SYNC_ARM",x,y)
  `define SET_DAC_COMMON_REG_CNTRL_1_EXT_SYNC_DISARM(x) SetField(DAC_COMMON_REG_CNTRL_1,"EXT_SYNC_DISARM",x)
  `define GET_DAC_COMMON_REG_CNTRL_1_EXT_SYNC_DISARM(x) GetField(DAC_COMMON_REG_CNTRL_1,"EXT_SYNC_DISARM",x)
  `define DEFAULT_DAC_COMMON_REG_CNTRL_1_EXT_SYNC_DISARM GetResetValue(DAC_COMMON_REG_CNTRL_1,"EXT_SYNC_DISARM")
  `define UPDATE_DAC_COMMON_REG_CNTRL_1_EXT_SYNC_DISARM(x,y) UpdateField(DAC_COMMON_REG_CNTRL_1,"EXT_SYNC_DISARM",x,y)
  `define SET_DAC_COMMON_REG_CNTRL_1_MANUAL_SYNC_REQUEST(x) SetField(DAC_COMMON_REG_CNTRL_1,"MANUAL_SYNC_REQUEST",x)
  `define GET_DAC_COMMON_REG_CNTRL_1_MANUAL_SYNC_REQUEST(x) GetField(DAC_COMMON_REG_CNTRL_1,"MANUAL_SYNC_REQUEST",x)
  `define DEFAULT_DAC_COMMON_REG_CNTRL_1_MANUAL_SYNC_REQUEST GetResetValue(DAC_COMMON_REG_CNTRL_1,"MANUAL_SYNC_REQUEST")
  `define UPDATE_DAC_COMMON_REG_CNTRL_1_MANUAL_SYNC_REQUEST(x,y) UpdateField(DAC_COMMON_REG_CNTRL_1,"MANUAL_SYNC_REQUEST",x,y)

  const reg_t DAC_COMMON_REG_CNTRL_2 = '{ 'h0048, "REG_CNTRL_2" , '{
    "SDR_DDR_N": '{ 16, 16, RW, 'h0 },
    "SYMB_OP": '{ 15, 15, RW, 'h0 },
    "SYMB_8_16B": '{ 14, 14, RW, 'h0 },
    "NUM_LANES": '{ 12, 8, RW, 'h0 },
    "PAR_TYPE": '{ 7, 7, RW, 'h0 },
    "PAR_ENB": '{ 6, 6, RW, 'h0 },
    "R1_MODE": '{ 5, 5, RW, 'h0 },
    "DATA_FORMAT": '{ 4, 4, RW, 'h0 }}};
  `define SET_DAC_COMMON_REG_CNTRL_2_SDR_DDR_N(x) SetField(DAC_COMMON_REG_CNTRL_2,"SDR_DDR_N",x)
  `define GET_DAC_COMMON_REG_CNTRL_2_SDR_DDR_N(x) GetField(DAC_COMMON_REG_CNTRL_2,"SDR_DDR_N",x)
  `define DEFAULT_DAC_COMMON_REG_CNTRL_2_SDR_DDR_N GetResetValue(DAC_COMMON_REG_CNTRL_2,"SDR_DDR_N")
  `define UPDATE_DAC_COMMON_REG_CNTRL_2_SDR_DDR_N(x,y) UpdateField(DAC_COMMON_REG_CNTRL_2,"SDR_DDR_N",x,y)
  `define SET_DAC_COMMON_REG_CNTRL_2_SYMB_OP(x) SetField(DAC_COMMON_REG_CNTRL_2,"SYMB_OP",x)
  `define GET_DAC_COMMON_REG_CNTRL_2_SYMB_OP(x) GetField(DAC_COMMON_REG_CNTRL_2,"SYMB_OP",x)
  `define DEFAULT_DAC_COMMON_REG_CNTRL_2_SYMB_OP GetResetValue(DAC_COMMON_REG_CNTRL_2,"SYMB_OP")
  `define UPDATE_DAC_COMMON_REG_CNTRL_2_SYMB_OP(x,y) UpdateField(DAC_COMMON_REG_CNTRL_2,"SYMB_OP",x,y)
  `define SET_DAC_COMMON_REG_CNTRL_2_SYMB_8_16B(x) SetField(DAC_COMMON_REG_CNTRL_2,"SYMB_8_16B",x)
  `define GET_DAC_COMMON_REG_CNTRL_2_SYMB_8_16B(x) GetField(DAC_COMMON_REG_CNTRL_2,"SYMB_8_16B",x)
  `define DEFAULT_DAC_COMMON_REG_CNTRL_2_SYMB_8_16B GetResetValue(DAC_COMMON_REG_CNTRL_2,"SYMB_8_16B")
  `define UPDATE_DAC_COMMON_REG_CNTRL_2_SYMB_8_16B(x,y) UpdateField(DAC_COMMON_REG_CNTRL_2,"SYMB_8_16B",x,y)
  `define SET_DAC_COMMON_REG_CNTRL_2_NUM_LANES(x) SetField(DAC_COMMON_REG_CNTRL_2,"NUM_LANES",x)
  `define GET_DAC_COMMON_REG_CNTRL_2_NUM_LANES(x) GetField(DAC_COMMON_REG_CNTRL_2,"NUM_LANES",x)
  `define DEFAULT_DAC_COMMON_REG_CNTRL_2_NUM_LANES GetResetValue(DAC_COMMON_REG_CNTRL_2,"NUM_LANES")
  `define UPDATE_DAC_COMMON_REG_CNTRL_2_NUM_LANES(x,y) UpdateField(DAC_COMMON_REG_CNTRL_2,"NUM_LANES",x,y)
  `define SET_DAC_COMMON_REG_CNTRL_2_PAR_TYPE(x) SetField(DAC_COMMON_REG_CNTRL_2,"PAR_TYPE",x)
  `define GET_DAC_COMMON_REG_CNTRL_2_PAR_TYPE(x) GetField(DAC_COMMON_REG_CNTRL_2,"PAR_TYPE",x)
  `define DEFAULT_DAC_COMMON_REG_CNTRL_2_PAR_TYPE GetResetValue(DAC_COMMON_REG_CNTRL_2,"PAR_TYPE")
  `define UPDATE_DAC_COMMON_REG_CNTRL_2_PAR_TYPE(x,y) UpdateField(DAC_COMMON_REG_CNTRL_2,"PAR_TYPE",x,y)
  `define SET_DAC_COMMON_REG_CNTRL_2_PAR_ENB(x) SetField(DAC_COMMON_REG_CNTRL_2,"PAR_ENB",x)
  `define GET_DAC_COMMON_REG_CNTRL_2_PAR_ENB(x) GetField(DAC_COMMON_REG_CNTRL_2,"PAR_ENB",x)
  `define DEFAULT_DAC_COMMON_REG_CNTRL_2_PAR_ENB GetResetValue(DAC_COMMON_REG_CNTRL_2,"PAR_ENB")
  `define UPDATE_DAC_COMMON_REG_CNTRL_2_PAR_ENB(x,y) UpdateField(DAC_COMMON_REG_CNTRL_2,"PAR_ENB",x,y)
  `define SET_DAC_COMMON_REG_CNTRL_2_R1_MODE(x) SetField(DAC_COMMON_REG_CNTRL_2,"R1_MODE",x)
  `define GET_DAC_COMMON_REG_CNTRL_2_R1_MODE(x) GetField(DAC_COMMON_REG_CNTRL_2,"R1_MODE",x)
  `define DEFAULT_DAC_COMMON_REG_CNTRL_2_R1_MODE GetResetValue(DAC_COMMON_REG_CNTRL_2,"R1_MODE")
  `define UPDATE_DAC_COMMON_REG_CNTRL_2_R1_MODE(x,y) UpdateField(DAC_COMMON_REG_CNTRL_2,"R1_MODE",x,y)
  `define SET_DAC_COMMON_REG_CNTRL_2_DATA_FORMAT(x) SetField(DAC_COMMON_REG_CNTRL_2,"DATA_FORMAT",x)
  `define GET_DAC_COMMON_REG_CNTRL_2_DATA_FORMAT(x) GetField(DAC_COMMON_REG_CNTRL_2,"DATA_FORMAT",x)
  `define DEFAULT_DAC_COMMON_REG_CNTRL_2_DATA_FORMAT GetResetValue(DAC_COMMON_REG_CNTRL_2,"DATA_FORMAT")
  `define UPDATE_DAC_COMMON_REG_CNTRL_2_DATA_FORMAT(x,y) UpdateField(DAC_COMMON_REG_CNTRL_2,"DATA_FORMAT",x,y)

  const reg_t DAC_COMMON_REG_RATECNTRL = '{ 'h004c, "REG_RATECNTRL" , '{
    "RATE": '{ 7, 0, RW, 'h00 }}};
  `define SET_DAC_COMMON_REG_RATECNTRL_RATE(x) SetField(DAC_COMMON_REG_RATECNTRL,"RATE",x)
  `define GET_DAC_COMMON_REG_RATECNTRL_RATE(x) GetField(DAC_COMMON_REG_RATECNTRL,"RATE",x)
  `define DEFAULT_DAC_COMMON_REG_RATECNTRL_RATE GetResetValue(DAC_COMMON_REG_RATECNTRL,"RATE")
  `define UPDATE_DAC_COMMON_REG_RATECNTRL_RATE(x,y) UpdateField(DAC_COMMON_REG_RATECNTRL,"RATE",x,y)

  const reg_t DAC_COMMON_REG_FRAME = '{ 'h0050, "REG_FRAME" , '{
    "FRAME": '{ 0, 0, RW, 'h0 }}};
  `define SET_DAC_COMMON_REG_FRAME_FRAME(x) SetField(DAC_COMMON_REG_FRAME,"FRAME",x)
  `define GET_DAC_COMMON_REG_FRAME_FRAME(x) GetField(DAC_COMMON_REG_FRAME,"FRAME",x)
  `define DEFAULT_DAC_COMMON_REG_FRAME_FRAME GetResetValue(DAC_COMMON_REG_FRAME,"FRAME")
  `define UPDATE_DAC_COMMON_REG_FRAME_FRAME(x,y) UpdateField(DAC_COMMON_REG_FRAME,"FRAME",x,y)

  const reg_t DAC_COMMON_REG_STATUS1 = '{ 'h0054, "REG_STATUS1" , '{
    "CLK_FREQ": '{ 31, 0, RO, 'h00000000 }}};
  `define SET_DAC_COMMON_REG_STATUS1_CLK_FREQ(x) SetField(DAC_COMMON_REG_STATUS1,"CLK_FREQ",x)
  `define GET_DAC_COMMON_REG_STATUS1_CLK_FREQ(x) GetField(DAC_COMMON_REG_STATUS1,"CLK_FREQ",x)
  `define DEFAULT_DAC_COMMON_REG_STATUS1_CLK_FREQ GetResetValue(DAC_COMMON_REG_STATUS1,"CLK_FREQ")
  `define UPDATE_DAC_COMMON_REG_STATUS1_CLK_FREQ(x,y) UpdateField(DAC_COMMON_REG_STATUS1,"CLK_FREQ",x,y)

  const reg_t DAC_COMMON_REG_STATUS2 = '{ 'h0058, "REG_STATUS2" , '{
    "CLK_RATIO": '{ 31, 0, RO, 'h00000000 }}};
  `define SET_DAC_COMMON_REG_STATUS2_CLK_RATIO(x) SetField(DAC_COMMON_REG_STATUS2,"CLK_RATIO",x)
  `define GET_DAC_COMMON_REG_STATUS2_CLK_RATIO(x) GetField(DAC_COMMON_REG_STATUS2,"CLK_RATIO",x)
  `define DEFAULT_DAC_COMMON_REG_STATUS2_CLK_RATIO GetResetValue(DAC_COMMON_REG_STATUS2,"CLK_RATIO")
  `define UPDATE_DAC_COMMON_REG_STATUS2_CLK_RATIO(x,y) UpdateField(DAC_COMMON_REG_STATUS2,"CLK_RATIO",x,y)

  const reg_t DAC_COMMON_REG_STATUS3 = '{ 'h005c, "REG_STATUS3" , '{
    "STATUS": '{ 0, 0, RO, 'h0 }}};
  `define SET_DAC_COMMON_REG_STATUS3_STATUS(x) SetField(DAC_COMMON_REG_STATUS3,"STATUS",x)
  `define GET_DAC_COMMON_REG_STATUS3_STATUS(x) GetField(DAC_COMMON_REG_STATUS3,"STATUS",x)
  `define DEFAULT_DAC_COMMON_REG_STATUS3_STATUS GetResetValue(DAC_COMMON_REG_STATUS3,"STATUS")
  `define UPDATE_DAC_COMMON_REG_STATUS3_STATUS(x,y) UpdateField(DAC_COMMON_REG_STATUS3,"STATUS",x,y)

  const reg_t DAC_COMMON_REG_DAC_CLKSEL = '{ 'h0060, "REG_DAC_CLKSEL" , '{
    "DAC_CLKSEL": '{ 0, 0, RW, 'h0 }}};
  `define SET_DAC_COMMON_REG_DAC_CLKSEL_DAC_CLKSEL(x) SetField(DAC_COMMON_REG_DAC_CLKSEL,"DAC_CLKSEL",x)
  `define GET_DAC_COMMON_REG_DAC_CLKSEL_DAC_CLKSEL(x) GetField(DAC_COMMON_REG_DAC_CLKSEL,"DAC_CLKSEL",x)
  `define DEFAULT_DAC_COMMON_REG_DAC_CLKSEL_DAC_CLKSEL GetResetValue(DAC_COMMON_REG_DAC_CLKSEL,"DAC_CLKSEL")
  `define UPDATE_DAC_COMMON_REG_DAC_CLKSEL_DAC_CLKSEL(x,y) UpdateField(DAC_COMMON_REG_DAC_CLKSEL,"DAC_CLKSEL",x,y)

  const reg_t DAC_COMMON_REG_SYNC_STATUS = '{ 'h0068, "REG_SYNC_STATUS" , '{
    "DAC_SYNC_STATUS": '{ 0, 0, RO, 'h0 }}};
  `define SET_DAC_COMMON_REG_SYNC_STATUS_DAC_SYNC_STATUS(x) SetField(DAC_COMMON_REG_SYNC_STATUS,"DAC_SYNC_STATUS",x)
  `define GET_DAC_COMMON_REG_SYNC_STATUS_DAC_SYNC_STATUS(x) GetField(DAC_COMMON_REG_SYNC_STATUS,"DAC_SYNC_STATUS",x)
  `define DEFAULT_DAC_COMMON_REG_SYNC_STATUS_DAC_SYNC_STATUS GetResetValue(DAC_COMMON_REG_SYNC_STATUS,"DAC_SYNC_STATUS")
  `define UPDATE_DAC_COMMON_REG_SYNC_STATUS_DAC_SYNC_STATUS(x,y) UpdateField(DAC_COMMON_REG_SYNC_STATUS,"DAC_SYNC_STATUS",x,y)

  const reg_t DAC_COMMON_REG_DRP_CNTRL = '{ 'h0070, "REG_DRP_CNTRL" , '{
    "DRP_RWN": '{ 28, 28, RW, 'h0 },
    "DRP_ADDRESS": '{ 27, 16, RW, 'h00 }}};
  `define SET_DAC_COMMON_REG_DRP_CNTRL_DRP_RWN(x) SetField(DAC_COMMON_REG_DRP_CNTRL,"DRP_RWN",x)
  `define GET_DAC_COMMON_REG_DRP_CNTRL_DRP_RWN(x) GetField(DAC_COMMON_REG_DRP_CNTRL,"DRP_RWN",x)
  `define DEFAULT_DAC_COMMON_REG_DRP_CNTRL_DRP_RWN GetResetValue(DAC_COMMON_REG_DRP_CNTRL,"DRP_RWN")
  `define UPDATE_DAC_COMMON_REG_DRP_CNTRL_DRP_RWN(x,y) UpdateField(DAC_COMMON_REG_DRP_CNTRL,"DRP_RWN",x,y)
  `define SET_DAC_COMMON_REG_DRP_CNTRL_DRP_ADDRESS(x) SetField(DAC_COMMON_REG_DRP_CNTRL,"DRP_ADDRESS",x)
  `define GET_DAC_COMMON_REG_DRP_CNTRL_DRP_ADDRESS(x) GetField(DAC_COMMON_REG_DRP_CNTRL,"DRP_ADDRESS",x)
  `define DEFAULT_DAC_COMMON_REG_DRP_CNTRL_DRP_ADDRESS GetResetValue(DAC_COMMON_REG_DRP_CNTRL,"DRP_ADDRESS")
  `define UPDATE_DAC_COMMON_REG_DRP_CNTRL_DRP_ADDRESS(x,y) UpdateField(DAC_COMMON_REG_DRP_CNTRL,"DRP_ADDRESS",x,y)

  const reg_t DAC_COMMON_REG_DRP_STATUS = '{ 'h0074, "REG_DRP_STATUS" , '{
    "DRP_LOCKED": '{ 17, 17, RO, 'h0 },
    "DRP_STATUS": '{ 16, 16, RO, 'h0 }}};
  `define SET_DAC_COMMON_REG_DRP_STATUS_DRP_LOCKED(x) SetField(DAC_COMMON_REG_DRP_STATUS,"DRP_LOCKED",x)
  `define GET_DAC_COMMON_REG_DRP_STATUS_DRP_LOCKED(x) GetField(DAC_COMMON_REG_DRP_STATUS,"DRP_LOCKED",x)
  `define DEFAULT_DAC_COMMON_REG_DRP_STATUS_DRP_LOCKED GetResetValue(DAC_COMMON_REG_DRP_STATUS,"DRP_LOCKED")
  `define UPDATE_DAC_COMMON_REG_DRP_STATUS_DRP_LOCKED(x,y) UpdateField(DAC_COMMON_REG_DRP_STATUS,"DRP_LOCKED",x,y)
  `define SET_DAC_COMMON_REG_DRP_STATUS_DRP_STATUS(x) SetField(DAC_COMMON_REG_DRP_STATUS,"DRP_STATUS",x)
  `define GET_DAC_COMMON_REG_DRP_STATUS_DRP_STATUS(x) GetField(DAC_COMMON_REG_DRP_STATUS,"DRP_STATUS",x)
  `define DEFAULT_DAC_COMMON_REG_DRP_STATUS_DRP_STATUS GetResetValue(DAC_COMMON_REG_DRP_STATUS,"DRP_STATUS")
  `define UPDATE_DAC_COMMON_REG_DRP_STATUS_DRP_STATUS(x,y) UpdateField(DAC_COMMON_REG_DRP_STATUS,"DRP_STATUS",x,y)

  const reg_t DAC_COMMON_REG_DRP_WDATA = '{ 'h0078, "REG_DRP_WDATA" , '{
    "DRP_WDATA": '{ 15, 0, RW, 'h0000 }}};
  `define SET_DAC_COMMON_REG_DRP_WDATA_DRP_WDATA(x) SetField(DAC_COMMON_REG_DRP_WDATA,"DRP_WDATA",x)
  `define GET_DAC_COMMON_REG_DRP_WDATA_DRP_WDATA(x) GetField(DAC_COMMON_REG_DRP_WDATA,"DRP_WDATA",x)
  `define DEFAULT_DAC_COMMON_REG_DRP_WDATA_DRP_WDATA GetResetValue(DAC_COMMON_REG_DRP_WDATA,"DRP_WDATA")
  `define UPDATE_DAC_COMMON_REG_DRP_WDATA_DRP_WDATA(x,y) UpdateField(DAC_COMMON_REG_DRP_WDATA,"DRP_WDATA",x,y)

  const reg_t DAC_COMMON_REG_DRP_RDATA = '{ 'h007c, "REG_DRP_RDATA" , '{
    "DRP_RDATA": '{ 15, 0, RO, 'h0000 }}};
  `define SET_DAC_COMMON_REG_DRP_RDATA_DRP_RDATA(x) SetField(DAC_COMMON_REG_DRP_RDATA,"DRP_RDATA",x)
  `define GET_DAC_COMMON_REG_DRP_RDATA_DRP_RDATA(x) GetField(DAC_COMMON_REG_DRP_RDATA,"DRP_RDATA",x)
  `define DEFAULT_DAC_COMMON_REG_DRP_RDATA_DRP_RDATA GetResetValue(DAC_COMMON_REG_DRP_RDATA,"DRP_RDATA")
  `define UPDATE_DAC_COMMON_REG_DRP_RDATA_DRP_RDATA(x,y) UpdateField(DAC_COMMON_REG_DRP_RDATA,"DRP_RDATA",x,y)

  const reg_t DAC_COMMON_REG_DAC_CUSTOM_RD = '{ 'h0080, "REG_DAC_CUSTOM_RD" , '{
    "DAC_CUSTOM_RD": '{ 31, 0, RO, 'h00000000 }}};
  `define SET_DAC_COMMON_REG_DAC_CUSTOM_RD_DAC_CUSTOM_RD(x) SetField(DAC_COMMON_REG_DAC_CUSTOM_RD,"DAC_CUSTOM_RD",x)
  `define GET_DAC_COMMON_REG_DAC_CUSTOM_RD_DAC_CUSTOM_RD(x) GetField(DAC_COMMON_REG_DAC_CUSTOM_RD,"DAC_CUSTOM_RD",x)
  `define DEFAULT_DAC_COMMON_REG_DAC_CUSTOM_RD_DAC_CUSTOM_RD GetResetValue(DAC_COMMON_REG_DAC_CUSTOM_RD,"DAC_CUSTOM_RD")
  `define UPDATE_DAC_COMMON_REG_DAC_CUSTOM_RD_DAC_CUSTOM_RD(x,y) UpdateField(DAC_COMMON_REG_DAC_CUSTOM_RD,"DAC_CUSTOM_RD",x,y)

  const reg_t DAC_COMMON_REG_DAC_CUSTOM_WR = '{ 'h0084, "REG_DAC_CUSTOM_WR" , '{
    "DAC_CUSTOM_WR": '{ 31, 0, RW, 'h00000000 }}};
  `define SET_DAC_COMMON_REG_DAC_CUSTOM_WR_DAC_CUSTOM_WR(x) SetField(DAC_COMMON_REG_DAC_CUSTOM_WR,"DAC_CUSTOM_WR",x)
  `define GET_DAC_COMMON_REG_DAC_CUSTOM_WR_DAC_CUSTOM_WR(x) GetField(DAC_COMMON_REG_DAC_CUSTOM_WR,"DAC_CUSTOM_WR",x)
  `define DEFAULT_DAC_COMMON_REG_DAC_CUSTOM_WR_DAC_CUSTOM_WR GetResetValue(DAC_COMMON_REG_DAC_CUSTOM_WR,"DAC_CUSTOM_WR")
  `define UPDATE_DAC_COMMON_REG_DAC_CUSTOM_WR_DAC_CUSTOM_WR(x,y) UpdateField(DAC_COMMON_REG_DAC_CUSTOM_WR,"DAC_CUSTOM_WR",x,y)

  const reg_t DAC_COMMON_REG_UI_STATUS = '{ 'h0088, "REG_UI_STATUS" , '{
    "IF_BUSY": '{ 4, 4, RO, 'h0 },
    "UI_OVF": '{ 1, 1, RW1C, 'h0 },
    "UI_UNF": '{ 0, 0, RW1C, 'h0 }}};
  `define SET_DAC_COMMON_REG_UI_STATUS_IF_BUSY(x) SetField(DAC_COMMON_REG_UI_STATUS,"IF_BUSY",x)
  `define GET_DAC_COMMON_REG_UI_STATUS_IF_BUSY(x) GetField(DAC_COMMON_REG_UI_STATUS,"IF_BUSY",x)
  `define DEFAULT_DAC_COMMON_REG_UI_STATUS_IF_BUSY GetResetValue(DAC_COMMON_REG_UI_STATUS,"IF_BUSY")
  `define UPDATE_DAC_COMMON_REG_UI_STATUS_IF_BUSY(x,y) UpdateField(DAC_COMMON_REG_UI_STATUS,"IF_BUSY",x,y)
  `define SET_DAC_COMMON_REG_UI_STATUS_UI_OVF(x) SetField(DAC_COMMON_REG_UI_STATUS,"UI_OVF",x)
  `define GET_DAC_COMMON_REG_UI_STATUS_UI_OVF(x) GetField(DAC_COMMON_REG_UI_STATUS,"UI_OVF",x)
  `define DEFAULT_DAC_COMMON_REG_UI_STATUS_UI_OVF GetResetValue(DAC_COMMON_REG_UI_STATUS,"UI_OVF")
  `define UPDATE_DAC_COMMON_REG_UI_STATUS_UI_OVF(x,y) UpdateField(DAC_COMMON_REG_UI_STATUS,"UI_OVF",x,y)
  `define SET_DAC_COMMON_REG_UI_STATUS_UI_UNF(x) SetField(DAC_COMMON_REG_UI_STATUS,"UI_UNF",x)
  `define GET_DAC_COMMON_REG_UI_STATUS_UI_UNF(x) GetField(DAC_COMMON_REG_UI_STATUS,"UI_UNF",x)
  `define DEFAULT_DAC_COMMON_REG_UI_STATUS_UI_UNF GetResetValue(DAC_COMMON_REG_UI_STATUS,"UI_UNF")
  `define UPDATE_DAC_COMMON_REG_UI_STATUS_UI_UNF(x,y) UpdateField(DAC_COMMON_REG_UI_STATUS,"UI_UNF",x,y)

  const reg_t DAC_COMMON_REG_DAC_CUSTOM_CTRL = '{ 'h008c, "REG_DAC_CUSTOM_CTRL" , '{
    "DAC_CUSTOM_CTRL": '{ 31, 0, RW, 'h00000000 }}};
  `define SET_DAC_COMMON_REG_DAC_CUSTOM_CTRL_DAC_CUSTOM_CTRL(x) SetField(DAC_COMMON_REG_DAC_CUSTOM_CTRL,"DAC_CUSTOM_CTRL",x)
  `define GET_DAC_COMMON_REG_DAC_CUSTOM_CTRL_DAC_CUSTOM_CTRL(x) GetField(DAC_COMMON_REG_DAC_CUSTOM_CTRL,"DAC_CUSTOM_CTRL",x)
  `define DEFAULT_DAC_COMMON_REG_DAC_CUSTOM_CTRL_DAC_CUSTOM_CTRL GetResetValue(DAC_COMMON_REG_DAC_CUSTOM_CTRL,"DAC_CUSTOM_CTRL")
  `define UPDATE_DAC_COMMON_REG_DAC_CUSTOM_CTRL_DAC_CUSTOM_CTRL(x,y) UpdateField(DAC_COMMON_REG_DAC_CUSTOM_CTRL,"DAC_CUSTOM_CTRL",x,y)

  const reg_t DAC_COMMON_REG_USR_CNTRL_1 = '{ 'h00a0, "REG_USR_CNTRL_1" , '{
    "USR_CHANMAX": '{ 7, 0, RW, 'h00 }}};
  `define SET_DAC_COMMON_REG_USR_CNTRL_1_USR_CHANMAX(x) SetField(DAC_COMMON_REG_USR_CNTRL_1,"USR_CHANMAX",x)
  `define GET_DAC_COMMON_REG_USR_CNTRL_1_USR_CHANMAX(x) GetField(DAC_COMMON_REG_USR_CNTRL_1,"USR_CHANMAX",x)
  `define DEFAULT_DAC_COMMON_REG_USR_CNTRL_1_USR_CHANMAX GetResetValue(DAC_COMMON_REG_USR_CNTRL_1,"USR_CHANMAX")
  `define UPDATE_DAC_COMMON_REG_USR_CNTRL_1_USR_CHANMAX(x,y) UpdateField(DAC_COMMON_REG_USR_CNTRL_1,"USR_CHANMAX",x,y)

  const reg_t DAC_COMMON_REG_DAC_GPIO_IN = '{ 'h00b8, "REG_DAC_GPIO_IN" , '{
    "DAC_GPIO_IN": '{ 31, 0, RO, 'h00000000 }}};
  `define SET_DAC_COMMON_REG_DAC_GPIO_IN_DAC_GPIO_IN(x) SetField(DAC_COMMON_REG_DAC_GPIO_IN,"DAC_GPIO_IN",x)
  `define GET_DAC_COMMON_REG_DAC_GPIO_IN_DAC_GPIO_IN(x) GetField(DAC_COMMON_REG_DAC_GPIO_IN,"DAC_GPIO_IN",x)
  `define DEFAULT_DAC_COMMON_REG_DAC_GPIO_IN_DAC_GPIO_IN GetResetValue(DAC_COMMON_REG_DAC_GPIO_IN,"DAC_GPIO_IN")
  `define UPDATE_DAC_COMMON_REG_DAC_GPIO_IN_DAC_GPIO_IN(x,y) UpdateField(DAC_COMMON_REG_DAC_GPIO_IN,"DAC_GPIO_IN",x,y)

  const reg_t DAC_COMMON_REG_DAC_GPIO_OUT = '{ 'h00bc, "REG_DAC_GPIO_OUT" , '{
    "DAC_GPIO_OUT": '{ 31, 0, RW, 'h00000000 }}};
  `define SET_DAC_COMMON_REG_DAC_GPIO_OUT_DAC_GPIO_OUT(x) SetField(DAC_COMMON_REG_DAC_GPIO_OUT,"DAC_GPIO_OUT",x)
  `define GET_DAC_COMMON_REG_DAC_GPIO_OUT_DAC_GPIO_OUT(x) GetField(DAC_COMMON_REG_DAC_GPIO_OUT,"DAC_GPIO_OUT",x)
  `define DEFAULT_DAC_COMMON_REG_DAC_GPIO_OUT_DAC_GPIO_OUT GetResetValue(DAC_COMMON_REG_DAC_GPIO_OUT,"DAC_GPIO_OUT")
  `define UPDATE_DAC_COMMON_REG_DAC_GPIO_OUT_DAC_GPIO_OUT(x,y) UpdateField(DAC_COMMON_REG_DAC_GPIO_OUT,"DAC_GPIO_OUT",x,y)


/* DAC Channel (axi_ad*) */

  const reg_t DAC_CHANNEL_REG_CHAN_CNTRL_1 = '{ 'h0400, "REG_CHAN_CNTRL_1" , '{
    "DDS_PHASE_DW": '{ 21, 16, R, 'h0000 },
    "DDS_SCALE_1": '{ 15, 0, RW, 'h0000 }}};
  `define SET_DAC_CHANNEL_REG_CHAN_CNTRL_1_DDS_PHASE_DW(x) SetField(DAC_CHANNEL_REG_CHAN_CNTRL_1,"DDS_PHASE_DW",x)
  `define GET_DAC_CHANNEL_REG_CHAN_CNTRL_1_DDS_PHASE_DW(x) GetField(DAC_CHANNEL_REG_CHAN_CNTRL_1,"DDS_PHASE_DW",x)
  `define DEFAULT_DAC_CHANNEL_REG_CHAN_CNTRL_1_DDS_PHASE_DW GetResetValue(DAC_CHANNEL_REG_CHAN_CNTRL_1,"DDS_PHASE_DW")
  `define UPDATE_DAC_CHANNEL_REG_CHAN_CNTRL_1_DDS_PHASE_DW(x,y) UpdateField(DAC_CHANNEL_REG_CHAN_CNTRL_1,"DDS_PHASE_DW",x,y)
  `define SET_DAC_CHANNEL_REG_CHAN_CNTRL_1_DDS_SCALE_1(x) SetField(DAC_CHANNEL_REG_CHAN_CNTRL_1,"DDS_SCALE_1",x)
  `define GET_DAC_CHANNEL_REG_CHAN_CNTRL_1_DDS_SCALE_1(x) GetField(DAC_CHANNEL_REG_CHAN_CNTRL_1,"DDS_SCALE_1",x)
  `define DEFAULT_DAC_CHANNEL_REG_CHAN_CNTRL_1_DDS_SCALE_1 GetResetValue(DAC_CHANNEL_REG_CHAN_CNTRL_1,"DDS_SCALE_1")
  `define UPDATE_DAC_CHANNEL_REG_CHAN_CNTRL_1_DDS_SCALE_1(x,y) UpdateField(DAC_CHANNEL_REG_CHAN_CNTRL_1,"DDS_SCALE_1",x,y)

  const reg_t DAC_CHANNEL_REG_CHAN_CNTRL_2 = '{ 'h0404, "REG_CHAN_CNTRL_2" , '{
    "DDS_INIT_1": '{ 31, 16, RW, 'h0000 },
    "DDS_INCR_1": '{ 15, 0, RW, 'h0000 }}};
  `define SET_DAC_CHANNEL_REG_CHAN_CNTRL_2_DDS_INIT_1(x) SetField(DAC_CHANNEL_REG_CHAN_CNTRL_2,"DDS_INIT_1",x)
  `define GET_DAC_CHANNEL_REG_CHAN_CNTRL_2_DDS_INIT_1(x) GetField(DAC_CHANNEL_REG_CHAN_CNTRL_2,"DDS_INIT_1",x)
  `define DEFAULT_DAC_CHANNEL_REG_CHAN_CNTRL_2_DDS_INIT_1 GetResetValue(DAC_CHANNEL_REG_CHAN_CNTRL_2,"DDS_INIT_1")
  `define UPDATE_DAC_CHANNEL_REG_CHAN_CNTRL_2_DDS_INIT_1(x,y) UpdateField(DAC_CHANNEL_REG_CHAN_CNTRL_2,"DDS_INIT_1",x,y)
  `define SET_DAC_CHANNEL_REG_CHAN_CNTRL_2_DDS_INCR_1(x) SetField(DAC_CHANNEL_REG_CHAN_CNTRL_2,"DDS_INCR_1",x)
  `define GET_DAC_CHANNEL_REG_CHAN_CNTRL_2_DDS_INCR_1(x) GetField(DAC_CHANNEL_REG_CHAN_CNTRL_2,"DDS_INCR_1",x)
  `define DEFAULT_DAC_CHANNEL_REG_CHAN_CNTRL_2_DDS_INCR_1 GetResetValue(DAC_CHANNEL_REG_CHAN_CNTRL_2,"DDS_INCR_1")
  `define UPDATE_DAC_CHANNEL_REG_CHAN_CNTRL_2_DDS_INCR_1(x,y) UpdateField(DAC_CHANNEL_REG_CHAN_CNTRL_2,"DDS_INCR_1",x,y)

  const reg_t DAC_CHANNEL_REG_CHAN_CNTRL_3 = '{ 'h0408, "REG_CHAN_CNTRL_3" , '{
    "DDS_SCALE_2": '{ 15, 0, RW, 'h0000 }}};
  `define SET_DAC_CHANNEL_REG_CHAN_CNTRL_3_DDS_SCALE_2(x) SetField(DAC_CHANNEL_REG_CHAN_CNTRL_3,"DDS_SCALE_2",x)
  `define GET_DAC_CHANNEL_REG_CHAN_CNTRL_3_DDS_SCALE_2(x) GetField(DAC_CHANNEL_REG_CHAN_CNTRL_3,"DDS_SCALE_2",x)
  `define DEFAULT_DAC_CHANNEL_REG_CHAN_CNTRL_3_DDS_SCALE_2 GetResetValue(DAC_CHANNEL_REG_CHAN_CNTRL_3,"DDS_SCALE_2")
  `define UPDATE_DAC_CHANNEL_REG_CHAN_CNTRL_3_DDS_SCALE_2(x,y) UpdateField(DAC_CHANNEL_REG_CHAN_CNTRL_3,"DDS_SCALE_2",x,y)

  const reg_t DAC_CHANNEL_REG_CHAN_CNTRL_4 = '{ 'h040c, "REG_CHAN_CNTRL_4" , '{
    "DDS_INIT_2": '{ 31, 16, RW, 'h0000 },
    "DDS_INCR_2": '{ 15, 0, RW, 'h0000 }}};
  `define SET_DAC_CHANNEL_REG_CHAN_CNTRL_4_DDS_INIT_2(x) SetField(DAC_CHANNEL_REG_CHAN_CNTRL_4,"DDS_INIT_2",x)
  `define GET_DAC_CHANNEL_REG_CHAN_CNTRL_4_DDS_INIT_2(x) GetField(DAC_CHANNEL_REG_CHAN_CNTRL_4,"DDS_INIT_2",x)
  `define DEFAULT_DAC_CHANNEL_REG_CHAN_CNTRL_4_DDS_INIT_2 GetResetValue(DAC_CHANNEL_REG_CHAN_CNTRL_4,"DDS_INIT_2")
  `define UPDATE_DAC_CHANNEL_REG_CHAN_CNTRL_4_DDS_INIT_2(x,y) UpdateField(DAC_CHANNEL_REG_CHAN_CNTRL_4,"DDS_INIT_2",x,y)
  `define SET_DAC_CHANNEL_REG_CHAN_CNTRL_4_DDS_INCR_2(x) SetField(DAC_CHANNEL_REG_CHAN_CNTRL_4,"DDS_INCR_2",x)
  `define GET_DAC_CHANNEL_REG_CHAN_CNTRL_4_DDS_INCR_2(x) GetField(DAC_CHANNEL_REG_CHAN_CNTRL_4,"DDS_INCR_2",x)
  `define DEFAULT_DAC_CHANNEL_REG_CHAN_CNTRL_4_DDS_INCR_2 GetResetValue(DAC_CHANNEL_REG_CHAN_CNTRL_4,"DDS_INCR_2")
  `define UPDATE_DAC_CHANNEL_REG_CHAN_CNTRL_4_DDS_INCR_2(x,y) UpdateField(DAC_CHANNEL_REG_CHAN_CNTRL_4,"DDS_INCR_2",x,y)

  const reg_t DAC_CHANNEL_REG_CHAN_CNTRL_5 = '{ 'h0410, "REG_CHAN_CNTRL_5" , '{
    "DDS_PATT_2": '{ 31, 16, RW, 'h0000 },
    "DDS_PATT_1": '{ 15, 0, RW, 'h0000 }}};
  `define SET_DAC_CHANNEL_REG_CHAN_CNTRL_5_DDS_PATT_2(x) SetField(DAC_CHANNEL_REG_CHAN_CNTRL_5,"DDS_PATT_2",x)
  `define GET_DAC_CHANNEL_REG_CHAN_CNTRL_5_DDS_PATT_2(x) GetField(DAC_CHANNEL_REG_CHAN_CNTRL_5,"DDS_PATT_2",x)
  `define DEFAULT_DAC_CHANNEL_REG_CHAN_CNTRL_5_DDS_PATT_2 GetResetValue(DAC_CHANNEL_REG_CHAN_CNTRL_5,"DDS_PATT_2")
  `define UPDATE_DAC_CHANNEL_REG_CHAN_CNTRL_5_DDS_PATT_2(x,y) UpdateField(DAC_CHANNEL_REG_CHAN_CNTRL_5,"DDS_PATT_2",x,y)
  `define SET_DAC_CHANNEL_REG_CHAN_CNTRL_5_DDS_PATT_1(x) SetField(DAC_CHANNEL_REG_CHAN_CNTRL_5,"DDS_PATT_1",x)
  `define GET_DAC_CHANNEL_REG_CHAN_CNTRL_5_DDS_PATT_1(x) GetField(DAC_CHANNEL_REG_CHAN_CNTRL_5,"DDS_PATT_1",x)
  `define DEFAULT_DAC_CHANNEL_REG_CHAN_CNTRL_5_DDS_PATT_1 GetResetValue(DAC_CHANNEL_REG_CHAN_CNTRL_5,"DDS_PATT_1")
  `define UPDATE_DAC_CHANNEL_REG_CHAN_CNTRL_5_DDS_PATT_1(x,y) UpdateField(DAC_CHANNEL_REG_CHAN_CNTRL_5,"DDS_PATT_1",x,y)

  const reg_t DAC_CHANNEL_REG_CHAN_CNTRL_6 = '{ 'h0414, "REG_CHAN_CNTRL_6" , '{
    "IQCOR_ENB": '{ 2, 2, RW, 'h0 },
    "DAC_LB_OWR": '{ 1, 1, RW, 'h0 },
    "DAC_PN_OWR": '{ 0, 0, RW, 'h0 }}};
  `define SET_DAC_CHANNEL_REG_CHAN_CNTRL_6_IQCOR_ENB(x) SetField(DAC_CHANNEL_REG_CHAN_CNTRL_6,"IQCOR_ENB",x)
  `define GET_DAC_CHANNEL_REG_CHAN_CNTRL_6_IQCOR_ENB(x) GetField(DAC_CHANNEL_REG_CHAN_CNTRL_6,"IQCOR_ENB",x)
  `define DEFAULT_DAC_CHANNEL_REG_CHAN_CNTRL_6_IQCOR_ENB GetResetValue(DAC_CHANNEL_REG_CHAN_CNTRL_6,"IQCOR_ENB")
  `define UPDATE_DAC_CHANNEL_REG_CHAN_CNTRL_6_IQCOR_ENB(x,y) UpdateField(DAC_CHANNEL_REG_CHAN_CNTRL_6,"IQCOR_ENB",x,y)
  `define SET_DAC_CHANNEL_REG_CHAN_CNTRL_6_DAC_LB_OWR(x) SetField(DAC_CHANNEL_REG_CHAN_CNTRL_6,"DAC_LB_OWR",x)
  `define GET_DAC_CHANNEL_REG_CHAN_CNTRL_6_DAC_LB_OWR(x) GetField(DAC_CHANNEL_REG_CHAN_CNTRL_6,"DAC_LB_OWR",x)
  `define DEFAULT_DAC_CHANNEL_REG_CHAN_CNTRL_6_DAC_LB_OWR GetResetValue(DAC_CHANNEL_REG_CHAN_CNTRL_6,"DAC_LB_OWR")
  `define UPDATE_DAC_CHANNEL_REG_CHAN_CNTRL_6_DAC_LB_OWR(x,y) UpdateField(DAC_CHANNEL_REG_CHAN_CNTRL_6,"DAC_LB_OWR",x,y)
  `define SET_DAC_CHANNEL_REG_CHAN_CNTRL_6_DAC_PN_OWR(x) SetField(DAC_CHANNEL_REG_CHAN_CNTRL_6,"DAC_PN_OWR",x)
  `define GET_DAC_CHANNEL_REG_CHAN_CNTRL_6_DAC_PN_OWR(x) GetField(DAC_CHANNEL_REG_CHAN_CNTRL_6,"DAC_PN_OWR",x)
  `define DEFAULT_DAC_CHANNEL_REG_CHAN_CNTRL_6_DAC_PN_OWR GetResetValue(DAC_CHANNEL_REG_CHAN_CNTRL_6,"DAC_PN_OWR")
  `define UPDATE_DAC_CHANNEL_REG_CHAN_CNTRL_6_DAC_PN_OWR(x,y) UpdateField(DAC_CHANNEL_REG_CHAN_CNTRL_6,"DAC_PN_OWR",x,y)

  const reg_t DAC_CHANNEL_REG_CHAN_CNTRL_7 = '{ 'h0418, "REG_CHAN_CNTRL_7" , '{
    "DAC_DDS_SEL": '{ 3, 0, RW, 'h00 }}};
  `define SET_DAC_CHANNEL_REG_CHAN_CNTRL_7_DAC_DDS_SEL(x) SetField(DAC_CHANNEL_REG_CHAN_CNTRL_7,"DAC_DDS_SEL",x)
  `define GET_DAC_CHANNEL_REG_CHAN_CNTRL_7_DAC_DDS_SEL(x) GetField(DAC_CHANNEL_REG_CHAN_CNTRL_7,"DAC_DDS_SEL",x)
  `define DEFAULT_DAC_CHANNEL_REG_CHAN_CNTRL_7_DAC_DDS_SEL GetResetValue(DAC_CHANNEL_REG_CHAN_CNTRL_7,"DAC_DDS_SEL")
  `define UPDATE_DAC_CHANNEL_REG_CHAN_CNTRL_7_DAC_DDS_SEL(x,y) UpdateField(DAC_CHANNEL_REG_CHAN_CNTRL_7,"DAC_DDS_SEL",x,y)

  const reg_t DAC_CHANNEL_REG_CHAN_CNTRL_8 = '{ 'h041c, "REG_CHAN_CNTRL_8" , '{
    "IQCOR_COEFF_1": '{ 31, 16, RW, 'h0000 },
    "IQCOR_COEFF_2": '{ 15, 0, RW, 'h0000 }}};
  `define SET_DAC_CHANNEL_REG_CHAN_CNTRL_8_IQCOR_COEFF_1(x) SetField(DAC_CHANNEL_REG_CHAN_CNTRL_8,"IQCOR_COEFF_1",x)
  `define GET_DAC_CHANNEL_REG_CHAN_CNTRL_8_IQCOR_COEFF_1(x) GetField(DAC_CHANNEL_REG_CHAN_CNTRL_8,"IQCOR_COEFF_1",x)
  `define DEFAULT_DAC_CHANNEL_REG_CHAN_CNTRL_8_IQCOR_COEFF_1 GetResetValue(DAC_CHANNEL_REG_CHAN_CNTRL_8,"IQCOR_COEFF_1")
  `define UPDATE_DAC_CHANNEL_REG_CHAN_CNTRL_8_IQCOR_COEFF_1(x,y) UpdateField(DAC_CHANNEL_REG_CHAN_CNTRL_8,"IQCOR_COEFF_1",x,y)
  `define SET_DAC_CHANNEL_REG_CHAN_CNTRL_8_IQCOR_COEFF_2(x) SetField(DAC_CHANNEL_REG_CHAN_CNTRL_8,"IQCOR_COEFF_2",x)
  `define GET_DAC_CHANNEL_REG_CHAN_CNTRL_8_IQCOR_COEFF_2(x) GetField(DAC_CHANNEL_REG_CHAN_CNTRL_8,"IQCOR_COEFF_2",x)
  `define DEFAULT_DAC_CHANNEL_REG_CHAN_CNTRL_8_IQCOR_COEFF_2 GetResetValue(DAC_CHANNEL_REG_CHAN_CNTRL_8,"IQCOR_COEFF_2")
  `define UPDATE_DAC_CHANNEL_REG_CHAN_CNTRL_8_IQCOR_COEFF_2(x,y) UpdateField(DAC_CHANNEL_REG_CHAN_CNTRL_8,"IQCOR_COEFF_2",x,y)

  const reg_t DAC_CHANNEL_REG_USR_CNTRL_3 = '{ 'h0420, "REG_USR_CNTRL_3" , '{
    "USR_DATATYPE_BE": '{ 25, 25, RW, 'h0 },
    "USR_DATATYPE_SIGNED": '{ 24, 24, RW, 'h0 },
    "USR_DATATYPE_SHIFT": '{ 23, 16, RW, 'h00 },
    "USR_DATATYPE_TOTAL_BITS": '{ 15, 8, RW, 'h00 },
    "USR_DATATYPE_BITS": '{ 7, 0, RW, 'h00 }}};
  `define SET_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_BE(x) SetField(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_BE",x)
  `define GET_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_BE(x) GetField(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_BE",x)
  `define DEFAULT_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_BE GetResetValue(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_BE")
  `define UPDATE_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_BE(x,y) UpdateField(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_BE",x,y)
  `define SET_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_SIGNED(x) SetField(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_SIGNED",x)
  `define GET_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_SIGNED(x) GetField(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_SIGNED",x)
  `define DEFAULT_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_SIGNED GetResetValue(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_SIGNED")
  `define UPDATE_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_SIGNED(x,y) UpdateField(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_SIGNED",x,y)
  `define SET_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_SHIFT(x) SetField(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_SHIFT",x)
  `define GET_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_SHIFT(x) GetField(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_SHIFT",x)
  `define DEFAULT_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_SHIFT GetResetValue(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_SHIFT")
  `define UPDATE_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_SHIFT(x,y) UpdateField(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_SHIFT",x,y)
  `define SET_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_TOTAL_BITS(x) SetField(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_TOTAL_BITS",x)
  `define GET_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_TOTAL_BITS(x) GetField(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_TOTAL_BITS",x)
  `define DEFAULT_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_TOTAL_BITS GetResetValue(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_TOTAL_BITS")
  `define UPDATE_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_TOTAL_BITS(x,y) UpdateField(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_TOTAL_BITS",x,y)
  `define SET_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_BITS(x) SetField(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_BITS",x)
  `define GET_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_BITS(x) GetField(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_BITS",x)
  `define DEFAULT_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_BITS GetResetValue(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_BITS")
  `define UPDATE_DAC_CHANNEL_REG_USR_CNTRL_3_USR_DATATYPE_BITS(x,y) UpdateField(DAC_CHANNEL_REG_USR_CNTRL_3,"USR_DATATYPE_BITS",x,y)

  const reg_t DAC_CHANNEL_REG_USR_CNTRL_4 = '{ 'h0424, "REG_USR_CNTRL_4" , '{
    "USR_INTERPOLATION_M": '{ 31, 16, RW, 'h0000 },
    "USR_INTERPOLATION_N": '{ 15, 0, RW, 'h0000 }}};
  `define SET_DAC_CHANNEL_REG_USR_CNTRL_4_USR_INTERPOLATION_M(x) SetField(DAC_CHANNEL_REG_USR_CNTRL_4,"USR_INTERPOLATION_M",x)
  `define GET_DAC_CHANNEL_REG_USR_CNTRL_4_USR_INTERPOLATION_M(x) GetField(DAC_CHANNEL_REG_USR_CNTRL_4,"USR_INTERPOLATION_M",x)
  `define DEFAULT_DAC_CHANNEL_REG_USR_CNTRL_4_USR_INTERPOLATION_M GetResetValue(DAC_CHANNEL_REG_USR_CNTRL_4,"USR_INTERPOLATION_M")
  `define UPDATE_DAC_CHANNEL_REG_USR_CNTRL_4_USR_INTERPOLATION_M(x,y) UpdateField(DAC_CHANNEL_REG_USR_CNTRL_4,"USR_INTERPOLATION_M",x,y)
  `define SET_DAC_CHANNEL_REG_USR_CNTRL_4_USR_INTERPOLATION_N(x) SetField(DAC_CHANNEL_REG_USR_CNTRL_4,"USR_INTERPOLATION_N",x)
  `define GET_DAC_CHANNEL_REG_USR_CNTRL_4_USR_INTERPOLATION_N(x) GetField(DAC_CHANNEL_REG_USR_CNTRL_4,"USR_INTERPOLATION_N",x)
  `define DEFAULT_DAC_CHANNEL_REG_USR_CNTRL_4_USR_INTERPOLATION_N GetResetValue(DAC_CHANNEL_REG_USR_CNTRL_4,"USR_INTERPOLATION_N")
  `define UPDATE_DAC_CHANNEL_REG_USR_CNTRL_4_USR_INTERPOLATION_N(x,y) UpdateField(DAC_CHANNEL_REG_USR_CNTRL_4,"USR_INTERPOLATION_N",x,y)

  const reg_t DAC_CHANNEL_REG_USR_CNTRL_5 = '{ 'h0428, "REG_USR_CNTRL_5" , '{
    "DAC_IQ_MODE": '{ 0, 0, RW, 'h0 },
    "DAC_IQ_SWAP": '{ 1, 1, RW, 'h0 }}};
  `define SET_DAC_CHANNEL_REG_USR_CNTRL_5_DAC_IQ_MODE(x) SetField(DAC_CHANNEL_REG_USR_CNTRL_5,"DAC_IQ_MODE",x)
  `define GET_DAC_CHANNEL_REG_USR_CNTRL_5_DAC_IQ_MODE(x) GetField(DAC_CHANNEL_REG_USR_CNTRL_5,"DAC_IQ_MODE",x)
  `define DEFAULT_DAC_CHANNEL_REG_USR_CNTRL_5_DAC_IQ_MODE GetResetValue(DAC_CHANNEL_REG_USR_CNTRL_5,"DAC_IQ_MODE")
  `define UPDATE_DAC_CHANNEL_REG_USR_CNTRL_5_DAC_IQ_MODE(x,y) UpdateField(DAC_CHANNEL_REG_USR_CNTRL_5,"DAC_IQ_MODE",x,y)
  `define SET_DAC_CHANNEL_REG_USR_CNTRL_5_DAC_IQ_SWAP(x) SetField(DAC_CHANNEL_REG_USR_CNTRL_5,"DAC_IQ_SWAP",x)
  `define GET_DAC_CHANNEL_REG_USR_CNTRL_5_DAC_IQ_SWAP(x) GetField(DAC_CHANNEL_REG_USR_CNTRL_5,"DAC_IQ_SWAP",x)
  `define DEFAULT_DAC_CHANNEL_REG_USR_CNTRL_5_DAC_IQ_SWAP GetResetValue(DAC_CHANNEL_REG_USR_CNTRL_5,"DAC_IQ_SWAP")
  `define UPDATE_DAC_CHANNEL_REG_USR_CNTRL_5_DAC_IQ_SWAP(x,y) UpdateField(DAC_CHANNEL_REG_USR_CNTRL_5,"DAC_IQ_SWAP",x,y)

  const reg_t DAC_CHANNEL_REG_CHAN_CNTRL_9 = '{ 'h042c, "REG_CHAN_CNTRL_9" , '{
    "DDS_INIT_1_EXTENDED": '{ 31, 16, RW, 'h0000 },
    "DDS_INCR_1_EXTENDED": '{ 15, 0, RW, 'h0000 }}};
  `define SET_DAC_CHANNEL_REG_CHAN_CNTRL_9_DDS_INIT_1_EXTENDED(x) SetField(DAC_CHANNEL_REG_CHAN_CNTRL_9,"DDS_INIT_1_EXTENDED",x)
  `define GET_DAC_CHANNEL_REG_CHAN_CNTRL_9_DDS_INIT_1_EXTENDED(x) GetField(DAC_CHANNEL_REG_CHAN_CNTRL_9,"DDS_INIT_1_EXTENDED",x)
  `define DEFAULT_DAC_CHANNEL_REG_CHAN_CNTRL_9_DDS_INIT_1_EXTENDED GetResetValue(DAC_CHANNEL_REG_CHAN_CNTRL_9,"DDS_INIT_1_EXTENDED")
  `define UPDATE_DAC_CHANNEL_REG_CHAN_CNTRL_9_DDS_INIT_1_EXTENDED(x,y) UpdateField(DAC_CHANNEL_REG_CHAN_CNTRL_9,"DDS_INIT_1_EXTENDED",x,y)
  `define SET_DAC_CHANNEL_REG_CHAN_CNTRL_9_DDS_INCR_1_EXTENDED(x) SetField(DAC_CHANNEL_REG_CHAN_CNTRL_9,"DDS_INCR_1_EXTENDED",x)
  `define GET_DAC_CHANNEL_REG_CHAN_CNTRL_9_DDS_INCR_1_EXTENDED(x) GetField(DAC_CHANNEL_REG_CHAN_CNTRL_9,"DDS_INCR_1_EXTENDED",x)
  `define DEFAULT_DAC_CHANNEL_REG_CHAN_CNTRL_9_DDS_INCR_1_EXTENDED GetResetValue(DAC_CHANNEL_REG_CHAN_CNTRL_9,"DDS_INCR_1_EXTENDED")
  `define UPDATE_DAC_CHANNEL_REG_CHAN_CNTRL_9_DDS_INCR_1_EXTENDED(x,y) UpdateField(DAC_CHANNEL_REG_CHAN_CNTRL_9,"DDS_INCR_1_EXTENDED",x,y)

  const reg_t DAC_CHANNEL_REG_CHAN_CNTRL_10 = '{ 'h0430, "REG_CHAN_CNTRL_10" , '{
    "DDS_INIT_2_EXTENDED": '{ 31, 16, RW, 'h0000 },
    "DDS_INCR_2_EXTENDED": '{ 15, 0, RW, 'h0000 }}};
  `define SET_DAC_CHANNEL_REG_CHAN_CNTRL_10_DDS_INIT_2_EXTENDED(x) SetField(DAC_CHANNEL_REG_CHAN_CNTRL_10,"DDS_INIT_2_EXTENDED",x)
  `define GET_DAC_CHANNEL_REG_CHAN_CNTRL_10_DDS_INIT_2_EXTENDED(x) GetField(DAC_CHANNEL_REG_CHAN_CNTRL_10,"DDS_INIT_2_EXTENDED",x)
  `define DEFAULT_DAC_CHANNEL_REG_CHAN_CNTRL_10_DDS_INIT_2_EXTENDED GetResetValue(DAC_CHANNEL_REG_CHAN_CNTRL_10,"DDS_INIT_2_EXTENDED")
  `define UPDATE_DAC_CHANNEL_REG_CHAN_CNTRL_10_DDS_INIT_2_EXTENDED(x,y) UpdateField(DAC_CHANNEL_REG_CHAN_CNTRL_10,"DDS_INIT_2_EXTENDED",x,y)
  `define SET_DAC_CHANNEL_REG_CHAN_CNTRL_10_DDS_INCR_2_EXTENDED(x) SetField(DAC_CHANNEL_REG_CHAN_CNTRL_10,"DDS_INCR_2_EXTENDED",x)
  `define GET_DAC_CHANNEL_REG_CHAN_CNTRL_10_DDS_INCR_2_EXTENDED(x) GetField(DAC_CHANNEL_REG_CHAN_CNTRL_10,"DDS_INCR_2_EXTENDED",x)
  `define DEFAULT_DAC_CHANNEL_REG_CHAN_CNTRL_10_DDS_INCR_2_EXTENDED GetResetValue(DAC_CHANNEL_REG_CHAN_CNTRL_10,"DDS_INCR_2_EXTENDED")
  `define UPDATE_DAC_CHANNEL_REG_CHAN_CNTRL_10_DDS_INCR_2_EXTENDED(x,y) UpdateField(DAC_CHANNEL_REG_CHAN_CNTRL_10,"DDS_INCR_2_EXTENDED",x,y)


endpackage
