// ***************************************************************************
// ***************************************************************************
// Copyright (C) 2014-2024 Analog Devices, Inc. All rights reserved.
//
// In this HDL repository, there are many different and unique modules, consisting
// of various HDL (Verilog or VHDL) components. The individual modules are
// developed independently, and may be accompanied by separate and unique license
// terms.
//
// The user should read each of these license terms, and understand the
// freedoms and responsibilities that he or she has by using this source/core.
//
// This core is distributed in the hope that it will be useful, but WITHOUT ANY
// WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR
// A PARTICULAR PURPOSE.
//
// Redistribution and use of source or resulting binaries, with or without modification
// of this file, are permitted under one of the following two license terms:
//
//   1. The GNU General Public License version 2 as published by the
//      Free Software Foundation, which can be found in the top level directory
//      of this repository (LICENSE_GPL2), and also online at:
//      <https://www.gnu.org/licenses/old-licenses/gpl-2.0.html>
//
// OR
//
//   2. An ADI specific BSD license, which can be found in the top level directory
//      of this repository (LICENSE_ADIBSD), and also on-line at:
//      https://github.com/analogdevicesinc/hdl/blob/main/LICENSE_ADIBSD
//      This will allow to generate bit files and not release the source code,
//      as long as it attaches to an ADI device.
//
// ***************************************************************************
// ***************************************************************************
/* Auto generated Register Map */
/* Thu Mar 28 13:22:23 2024 */

package adi_regmap_fan_control_pkg;
  import adi_regmap_pkg::*;


/* Fan Controller (axi_fan_control) */

  const reg_t AXI_FAN_CONTROL_VERSION = '{ 'h0000, "VERSION" , '{
    "VERSION_MAJOR": '{ 31, 16, RO, 'h0001 },
    "VERSION_MINOR": '{ 15, 8, RO, 'h00 },
    "VERSION_PATCH": '{ 7, 0, RO, 'h61 }}};
  `define SET_AXI_FAN_CONTROL_VERSION_VERSION_MAJOR(x) SetField(AXI_FAN_CONTROL_VERSION,"VERSION_MAJOR",x)
  `define GET_AXI_FAN_CONTROL_VERSION_VERSION_MAJOR(x) GetField(AXI_FAN_CONTROL_VERSION,"VERSION_MAJOR",x)
  `define DEFAULT_AXI_FAN_CONTROL_VERSION_VERSION_MAJOR GetResetValue(AXI_FAN_CONTROL_VERSION,"VERSION_MAJOR")
  `define UPDATE_AXI_FAN_CONTROL_VERSION_VERSION_MAJOR(x,y) UpdateField(AXI_FAN_CONTROL_VERSION,"VERSION_MAJOR",x,y)
  `define SET_AXI_FAN_CONTROL_VERSION_VERSION_MINOR(x) SetField(AXI_FAN_CONTROL_VERSION,"VERSION_MINOR",x)
  `define GET_AXI_FAN_CONTROL_VERSION_VERSION_MINOR(x) GetField(AXI_FAN_CONTROL_VERSION,"VERSION_MINOR",x)
  `define DEFAULT_AXI_FAN_CONTROL_VERSION_VERSION_MINOR GetResetValue(AXI_FAN_CONTROL_VERSION,"VERSION_MINOR")
  `define UPDATE_AXI_FAN_CONTROL_VERSION_VERSION_MINOR(x,y) UpdateField(AXI_FAN_CONTROL_VERSION,"VERSION_MINOR",x,y)
  `define SET_AXI_FAN_CONTROL_VERSION_VERSION_PATCH(x) SetField(AXI_FAN_CONTROL_VERSION,"VERSION_PATCH",x)
  `define GET_AXI_FAN_CONTROL_VERSION_VERSION_PATCH(x) GetField(AXI_FAN_CONTROL_VERSION,"VERSION_PATCH",x)
  `define DEFAULT_AXI_FAN_CONTROL_VERSION_VERSION_PATCH GetResetValue(AXI_FAN_CONTROL_VERSION,"VERSION_PATCH")
  `define UPDATE_AXI_FAN_CONTROL_VERSION_VERSION_PATCH(x,y) UpdateField(AXI_FAN_CONTROL_VERSION,"VERSION_PATCH",x,y)

  const reg_t AXI_FAN_CONTROL_PERIPHERAL_ID = '{ 'h0004, "PERIPHERAL_ID" , '{
    "PERIPHERAL_ID": '{ 31, 0, RO, 0 }}};
  `define SET_AXI_FAN_CONTROL_PERIPHERAL_ID_PERIPHERAL_ID(x) SetField(AXI_FAN_CONTROL_PERIPHERAL_ID,"PERIPHERAL_ID",x)
  `define GET_AXI_FAN_CONTROL_PERIPHERAL_ID_PERIPHERAL_ID(x) GetField(AXI_FAN_CONTROL_PERIPHERAL_ID,"PERIPHERAL_ID",x)
  `define DEFAULT_AXI_FAN_CONTROL_PERIPHERAL_ID_PERIPHERAL_ID GetResetValue(AXI_FAN_CONTROL_PERIPHERAL_ID,"PERIPHERAL_ID")
  `define UPDATE_AXI_FAN_CONTROL_PERIPHERAL_ID_PERIPHERAL_ID(x,y) UpdateField(AXI_FAN_CONTROL_PERIPHERAL_ID,"PERIPHERAL_ID",x,y)

  const reg_t AXI_FAN_CONTROL_SCRATCH = '{ 'h0008, "SCRATCH" , '{
    "SCRATCH": '{ 31, 0, RW, 'h00000000 }}};
  `define SET_AXI_FAN_CONTROL_SCRATCH_SCRATCH(x) SetField(AXI_FAN_CONTROL_SCRATCH,"SCRATCH",x)
  `define GET_AXI_FAN_CONTROL_SCRATCH_SCRATCH(x) GetField(AXI_FAN_CONTROL_SCRATCH,"SCRATCH",x)
  `define DEFAULT_AXI_FAN_CONTROL_SCRATCH_SCRATCH GetResetValue(AXI_FAN_CONTROL_SCRATCH,"SCRATCH")
  `define UPDATE_AXI_FAN_CONTROL_SCRATCH_SCRATCH(x,y) UpdateField(AXI_FAN_CONTROL_SCRATCH,"SCRATCH",x,y)

  const reg_t AXI_FAN_CONTROL_IDENTIFICATION = '{ 'h000c, "IDENTIFICATION" , '{
    "IDENTIFICATION": '{ 31, 0, RO, 'h46414E43 }}};
  `define SET_AXI_FAN_CONTROL_IDENTIFICATION_IDENTIFICATION(x) SetField(AXI_FAN_CONTROL_IDENTIFICATION,"IDENTIFICATION",x)
  `define GET_AXI_FAN_CONTROL_IDENTIFICATION_IDENTIFICATION(x) GetField(AXI_FAN_CONTROL_IDENTIFICATION,"IDENTIFICATION",x)
  `define DEFAULT_AXI_FAN_CONTROL_IDENTIFICATION_IDENTIFICATION GetResetValue(AXI_FAN_CONTROL_IDENTIFICATION,"IDENTIFICATION")
  `define UPDATE_AXI_FAN_CONTROL_IDENTIFICATION_IDENTIFICATION(x,y) UpdateField(AXI_FAN_CONTROL_IDENTIFICATION,"IDENTIFICATION",x,y)

  const reg_t AXI_FAN_CONTROL_IRQ_MASK = '{ 'h0040, "IRQ_MASK" , '{
    "NEW_TACHO_MEASUREMENT": '{ 3, 3, RW, 'h1 },
    "TEMP_INCREASE": '{ 2, 2, RW, 'h1 },
    "TACHO_ERR": '{ 1, 1, RW, 'h1 },
    "PWM_CHANGED": '{ 0, 0, RW, 'h1 }}};
  `define SET_AXI_FAN_CONTROL_IRQ_MASK_NEW_TACHO_MEASUREMENT(x) SetField(AXI_FAN_CONTROL_IRQ_MASK,"NEW_TACHO_MEASUREMENT",x)
  `define GET_AXI_FAN_CONTROL_IRQ_MASK_NEW_TACHO_MEASUREMENT(x) GetField(AXI_FAN_CONTROL_IRQ_MASK,"NEW_TACHO_MEASUREMENT",x)
  `define DEFAULT_AXI_FAN_CONTROL_IRQ_MASK_NEW_TACHO_MEASUREMENT GetResetValue(AXI_FAN_CONTROL_IRQ_MASK,"NEW_TACHO_MEASUREMENT")
  `define UPDATE_AXI_FAN_CONTROL_IRQ_MASK_NEW_TACHO_MEASUREMENT(x,y) UpdateField(AXI_FAN_CONTROL_IRQ_MASK,"NEW_TACHO_MEASUREMENT",x,y)
  `define SET_AXI_FAN_CONTROL_IRQ_MASK_TEMP_INCREASE(x) SetField(AXI_FAN_CONTROL_IRQ_MASK,"TEMP_INCREASE",x)
  `define GET_AXI_FAN_CONTROL_IRQ_MASK_TEMP_INCREASE(x) GetField(AXI_FAN_CONTROL_IRQ_MASK,"TEMP_INCREASE",x)
  `define DEFAULT_AXI_FAN_CONTROL_IRQ_MASK_TEMP_INCREASE GetResetValue(AXI_FAN_CONTROL_IRQ_MASK,"TEMP_INCREASE")
  `define UPDATE_AXI_FAN_CONTROL_IRQ_MASK_TEMP_INCREASE(x,y) UpdateField(AXI_FAN_CONTROL_IRQ_MASK,"TEMP_INCREASE",x,y)
  `define SET_AXI_FAN_CONTROL_IRQ_MASK_TACHO_ERR(x) SetField(AXI_FAN_CONTROL_IRQ_MASK,"TACHO_ERR",x)
  `define GET_AXI_FAN_CONTROL_IRQ_MASK_TACHO_ERR(x) GetField(AXI_FAN_CONTROL_IRQ_MASK,"TACHO_ERR",x)
  `define DEFAULT_AXI_FAN_CONTROL_IRQ_MASK_TACHO_ERR GetResetValue(AXI_FAN_CONTROL_IRQ_MASK,"TACHO_ERR")
  `define UPDATE_AXI_FAN_CONTROL_IRQ_MASK_TACHO_ERR(x,y) UpdateField(AXI_FAN_CONTROL_IRQ_MASK,"TACHO_ERR",x,y)
  `define SET_AXI_FAN_CONTROL_IRQ_MASK_PWM_CHANGED(x) SetField(AXI_FAN_CONTROL_IRQ_MASK,"PWM_CHANGED",x)
  `define GET_AXI_FAN_CONTROL_IRQ_MASK_PWM_CHANGED(x) GetField(AXI_FAN_CONTROL_IRQ_MASK,"PWM_CHANGED",x)
  `define DEFAULT_AXI_FAN_CONTROL_IRQ_MASK_PWM_CHANGED GetResetValue(AXI_FAN_CONTROL_IRQ_MASK,"PWM_CHANGED")
  `define UPDATE_AXI_FAN_CONTROL_IRQ_MASK_PWM_CHANGED(x,y) UpdateField(AXI_FAN_CONTROL_IRQ_MASK,"PWM_CHANGED",x,y)

  const reg_t AXI_FAN_CONTROL_IRQ_PENDING = '{ 'h0044, "IRQ_PENDING" , '{
    "NEW_TACHO_MEASUREMENT": '{ 3, 3, RW1C, 'h0 },
    "TEMP_INCREASE": '{ 2, 2, RW1C, 'h0 },
    "TACHO_ERR": '{ 1, 1, RW1C, 'h0 },
    "PWM_CHANGED": '{ 0, 0, RW1C, 'h0 }}};
  `define SET_AXI_FAN_CONTROL_IRQ_PENDING_NEW_TACHO_MEASUREMENT(x) SetField(AXI_FAN_CONTROL_IRQ_PENDING,"NEW_TACHO_MEASUREMENT",x)
  `define GET_AXI_FAN_CONTROL_IRQ_PENDING_NEW_TACHO_MEASUREMENT(x) GetField(AXI_FAN_CONTROL_IRQ_PENDING,"NEW_TACHO_MEASUREMENT",x)
  `define DEFAULT_AXI_FAN_CONTROL_IRQ_PENDING_NEW_TACHO_MEASUREMENT GetResetValue(AXI_FAN_CONTROL_IRQ_PENDING,"NEW_TACHO_MEASUREMENT")
  `define UPDATE_AXI_FAN_CONTROL_IRQ_PENDING_NEW_TACHO_MEASUREMENT(x,y) UpdateField(AXI_FAN_CONTROL_IRQ_PENDING,"NEW_TACHO_MEASUREMENT",x,y)
  `define SET_AXI_FAN_CONTROL_IRQ_PENDING_TEMP_INCREASE(x) SetField(AXI_FAN_CONTROL_IRQ_PENDING,"TEMP_INCREASE",x)
  `define GET_AXI_FAN_CONTROL_IRQ_PENDING_TEMP_INCREASE(x) GetField(AXI_FAN_CONTROL_IRQ_PENDING,"TEMP_INCREASE",x)
  `define DEFAULT_AXI_FAN_CONTROL_IRQ_PENDING_TEMP_INCREASE GetResetValue(AXI_FAN_CONTROL_IRQ_PENDING,"TEMP_INCREASE")
  `define UPDATE_AXI_FAN_CONTROL_IRQ_PENDING_TEMP_INCREASE(x,y) UpdateField(AXI_FAN_CONTROL_IRQ_PENDING,"TEMP_INCREASE",x,y)
  `define SET_AXI_FAN_CONTROL_IRQ_PENDING_TACHO_ERR(x) SetField(AXI_FAN_CONTROL_IRQ_PENDING,"TACHO_ERR",x)
  `define GET_AXI_FAN_CONTROL_IRQ_PENDING_TACHO_ERR(x) GetField(AXI_FAN_CONTROL_IRQ_PENDING,"TACHO_ERR",x)
  `define DEFAULT_AXI_FAN_CONTROL_IRQ_PENDING_TACHO_ERR GetResetValue(AXI_FAN_CONTROL_IRQ_PENDING,"TACHO_ERR")
  `define UPDATE_AXI_FAN_CONTROL_IRQ_PENDING_TACHO_ERR(x,y) UpdateField(AXI_FAN_CONTROL_IRQ_PENDING,"TACHO_ERR",x,y)
  `define SET_AXI_FAN_CONTROL_IRQ_PENDING_PWM_CHANGED(x) SetField(AXI_FAN_CONTROL_IRQ_PENDING,"PWM_CHANGED",x)
  `define GET_AXI_FAN_CONTROL_IRQ_PENDING_PWM_CHANGED(x) GetField(AXI_FAN_CONTROL_IRQ_PENDING,"PWM_CHANGED",x)
  `define DEFAULT_AXI_FAN_CONTROL_IRQ_PENDING_PWM_CHANGED GetResetValue(AXI_FAN_CONTROL_IRQ_PENDING,"PWM_CHANGED")
  `define UPDATE_AXI_FAN_CONTROL_IRQ_PENDING_PWM_CHANGED(x,y) UpdateField(AXI_FAN_CONTROL_IRQ_PENDING,"PWM_CHANGED",x,y)

  const reg_t AXI_FAN_CONTROL_IRQ_SOURCE = '{ 'h0048, "IRQ_SOURCE" , '{
    "NEW_TACHO_MEASUREMENT": '{ 3, 3, RO, 'h0 },
    "TEMP_INCREASE": '{ 2, 2, RO, 'h0 },
    "TACHO_ERR": '{ 1, 1, RO, 'h0 },
    "PWM_CHANGED": '{ 0, 0, RO, 'h0 }}};
  `define SET_AXI_FAN_CONTROL_IRQ_SOURCE_NEW_TACHO_MEASUREMENT(x) SetField(AXI_FAN_CONTROL_IRQ_SOURCE,"NEW_TACHO_MEASUREMENT",x)
  `define GET_AXI_FAN_CONTROL_IRQ_SOURCE_NEW_TACHO_MEASUREMENT(x) GetField(AXI_FAN_CONTROL_IRQ_SOURCE,"NEW_TACHO_MEASUREMENT",x)
  `define DEFAULT_AXI_FAN_CONTROL_IRQ_SOURCE_NEW_TACHO_MEASUREMENT GetResetValue(AXI_FAN_CONTROL_IRQ_SOURCE,"NEW_TACHO_MEASUREMENT")
  `define UPDATE_AXI_FAN_CONTROL_IRQ_SOURCE_NEW_TACHO_MEASUREMENT(x,y) UpdateField(AXI_FAN_CONTROL_IRQ_SOURCE,"NEW_TACHO_MEASUREMENT",x,y)
  `define SET_AXI_FAN_CONTROL_IRQ_SOURCE_TEMP_INCREASE(x) SetField(AXI_FAN_CONTROL_IRQ_SOURCE,"TEMP_INCREASE",x)
  `define GET_AXI_FAN_CONTROL_IRQ_SOURCE_TEMP_INCREASE(x) GetField(AXI_FAN_CONTROL_IRQ_SOURCE,"TEMP_INCREASE",x)
  `define DEFAULT_AXI_FAN_CONTROL_IRQ_SOURCE_TEMP_INCREASE GetResetValue(AXI_FAN_CONTROL_IRQ_SOURCE,"TEMP_INCREASE")
  `define UPDATE_AXI_FAN_CONTROL_IRQ_SOURCE_TEMP_INCREASE(x,y) UpdateField(AXI_FAN_CONTROL_IRQ_SOURCE,"TEMP_INCREASE",x,y)
  `define SET_AXI_FAN_CONTROL_IRQ_SOURCE_TACHO_ERR(x) SetField(AXI_FAN_CONTROL_IRQ_SOURCE,"TACHO_ERR",x)
  `define GET_AXI_FAN_CONTROL_IRQ_SOURCE_TACHO_ERR(x) GetField(AXI_FAN_CONTROL_IRQ_SOURCE,"TACHO_ERR",x)
  `define DEFAULT_AXI_FAN_CONTROL_IRQ_SOURCE_TACHO_ERR GetResetValue(AXI_FAN_CONTROL_IRQ_SOURCE,"TACHO_ERR")
  `define UPDATE_AXI_FAN_CONTROL_IRQ_SOURCE_TACHO_ERR(x,y) UpdateField(AXI_FAN_CONTROL_IRQ_SOURCE,"TACHO_ERR",x,y)
  `define SET_AXI_FAN_CONTROL_IRQ_SOURCE_PWM_CHANGED(x) SetField(AXI_FAN_CONTROL_IRQ_SOURCE,"PWM_CHANGED",x)
  `define GET_AXI_FAN_CONTROL_IRQ_SOURCE_PWM_CHANGED(x) GetField(AXI_FAN_CONTROL_IRQ_SOURCE,"PWM_CHANGED",x)
  `define DEFAULT_AXI_FAN_CONTROL_IRQ_SOURCE_PWM_CHANGED GetResetValue(AXI_FAN_CONTROL_IRQ_SOURCE,"PWM_CHANGED")
  `define UPDATE_AXI_FAN_CONTROL_IRQ_SOURCE_PWM_CHANGED(x,y) UpdateField(AXI_FAN_CONTROL_IRQ_SOURCE,"PWM_CHANGED",x,y)

  const reg_t AXI_FAN_CONTROL_REG_RSTN = '{ 'h0080, "REG_RSTN" , '{
    "RSTN": '{ 0, 0, RW, 'h0 }}};
  `define SET_AXI_FAN_CONTROL_REG_RSTN_RSTN(x) SetField(AXI_FAN_CONTROL_REG_RSTN,"RSTN",x)
  `define GET_AXI_FAN_CONTROL_REG_RSTN_RSTN(x) GetField(AXI_FAN_CONTROL_REG_RSTN,"RSTN",x)
  `define DEFAULT_AXI_FAN_CONTROL_REG_RSTN_RSTN GetResetValue(AXI_FAN_CONTROL_REG_RSTN,"RSTN")
  `define UPDATE_AXI_FAN_CONTROL_REG_RSTN_RSTN(x,y) UpdateField(AXI_FAN_CONTROL_REG_RSTN,"RSTN",x,y)

  const reg_t AXI_FAN_CONTROL_PWM_WIDTH = '{ 'h0084, "PWM_WIDTH" , '{
    "PWM_WIDTH": '{ 31, 0, RW, 0 }}};
  `define SET_AXI_FAN_CONTROL_PWM_WIDTH_PWM_WIDTH(x) SetField(AXI_FAN_CONTROL_PWM_WIDTH,"PWM_WIDTH",x)
  `define GET_AXI_FAN_CONTROL_PWM_WIDTH_PWM_WIDTH(x) GetField(AXI_FAN_CONTROL_PWM_WIDTH,"PWM_WIDTH",x)
  `define DEFAULT_AXI_FAN_CONTROL_PWM_WIDTH_PWM_WIDTH GetResetValue(AXI_FAN_CONTROL_PWM_WIDTH,"PWM_WIDTH")
  `define UPDATE_AXI_FAN_CONTROL_PWM_WIDTH_PWM_WIDTH(x,y) UpdateField(AXI_FAN_CONTROL_PWM_WIDTH,"PWM_WIDTH",x,y)

  const reg_t AXI_FAN_CONTROL_TACHO_PERIOD = '{ 'h0088, "TACHO_PERIOD" , '{
    "TACHO_PERIOD": '{ 31, 0, RW, 'h00000000 }}};
  `define SET_AXI_FAN_CONTROL_TACHO_PERIOD_TACHO_PERIOD(x) SetField(AXI_FAN_CONTROL_TACHO_PERIOD,"TACHO_PERIOD",x)
  `define GET_AXI_FAN_CONTROL_TACHO_PERIOD_TACHO_PERIOD(x) GetField(AXI_FAN_CONTROL_TACHO_PERIOD,"TACHO_PERIOD",x)
  `define DEFAULT_AXI_FAN_CONTROL_TACHO_PERIOD_TACHO_PERIOD GetResetValue(AXI_FAN_CONTROL_TACHO_PERIOD,"TACHO_PERIOD")
  `define UPDATE_AXI_FAN_CONTROL_TACHO_PERIOD_TACHO_PERIOD(x,y) UpdateField(AXI_FAN_CONTROL_TACHO_PERIOD,"TACHO_PERIOD",x,y)

  const reg_t AXI_FAN_CONTROL_TACHO_TOLERANCE = '{ 'h008c, "TACHO_TOLERANCE" , '{
    "TACHO_TOLERANCE": '{ 31, 0, RW, 'h00000000 }}};
  `define SET_AXI_FAN_CONTROL_TACHO_TOLERANCE_TACHO_TOLERANCE(x) SetField(AXI_FAN_CONTROL_TACHO_TOLERANCE,"TACHO_TOLERANCE",x)
  `define GET_AXI_FAN_CONTROL_TACHO_TOLERANCE_TACHO_TOLERANCE(x) GetField(AXI_FAN_CONTROL_TACHO_TOLERANCE,"TACHO_TOLERANCE",x)
  `define DEFAULT_AXI_FAN_CONTROL_TACHO_TOLERANCE_TACHO_TOLERANCE GetResetValue(AXI_FAN_CONTROL_TACHO_TOLERANCE,"TACHO_TOLERANCE")
  `define UPDATE_AXI_FAN_CONTROL_TACHO_TOLERANCE_TACHO_TOLERANCE(x,y) UpdateField(AXI_FAN_CONTROL_TACHO_TOLERANCE,"TACHO_TOLERANCE",x,y)

  const reg_t AXI_FAN_CONTROL_TEMP_DATA_SOURCE = '{ 'h0090, "TEMP_DATA_SOURCE" , '{
    "TEMP_DATA_SOURCE": '{ 31, 0, RO, 0 }}};
  `define SET_AXI_FAN_CONTROL_TEMP_DATA_SOURCE_TEMP_DATA_SOURCE(x) SetField(AXI_FAN_CONTROL_TEMP_DATA_SOURCE,"TEMP_DATA_SOURCE",x)
  `define GET_AXI_FAN_CONTROL_TEMP_DATA_SOURCE_TEMP_DATA_SOURCE(x) GetField(AXI_FAN_CONTROL_TEMP_DATA_SOURCE,"TEMP_DATA_SOURCE",x)
  `define DEFAULT_AXI_FAN_CONTROL_TEMP_DATA_SOURCE_TEMP_DATA_SOURCE GetResetValue(AXI_FAN_CONTROL_TEMP_DATA_SOURCE,"TEMP_DATA_SOURCE")
  `define UPDATE_AXI_FAN_CONTROL_TEMP_DATA_SOURCE_TEMP_DATA_SOURCE(x,y) UpdateField(AXI_FAN_CONTROL_TEMP_DATA_SOURCE,"TEMP_DATA_SOURCE",x,y)

  const reg_t AXI_FAN_CONTROL_PWM_PERIOD = '{ 'h00c0, "PWM_PERIOD" , '{
    "PWM_PERIOD": '{ 31, 0, RO, 'h4E20 }}};
  `define SET_AXI_FAN_CONTROL_PWM_PERIOD_PWM_PERIOD(x) SetField(AXI_FAN_CONTROL_PWM_PERIOD,"PWM_PERIOD",x)
  `define GET_AXI_FAN_CONTROL_PWM_PERIOD_PWM_PERIOD(x) GetField(AXI_FAN_CONTROL_PWM_PERIOD,"PWM_PERIOD",x)
  `define DEFAULT_AXI_FAN_CONTROL_PWM_PERIOD_PWM_PERIOD GetResetValue(AXI_FAN_CONTROL_PWM_PERIOD,"PWM_PERIOD")
  `define UPDATE_AXI_FAN_CONTROL_PWM_PERIOD_PWM_PERIOD(x,y) UpdateField(AXI_FAN_CONTROL_PWM_PERIOD,"PWM_PERIOD",x,y)

  const reg_t AXI_FAN_CONTROL_TACHO_MEASUREMENT = '{ 'h00c4, "TACHO_MEASUREMENT" , '{
    "TACHO_MEASUREMENT": '{ 31, 0, RO, 'h00000000 }}};
  `define SET_AXI_FAN_CONTROL_TACHO_MEASUREMENT_TACHO_MEASUREMENT(x) SetField(AXI_FAN_CONTROL_TACHO_MEASUREMENT,"TACHO_MEASUREMENT",x)
  `define GET_AXI_FAN_CONTROL_TACHO_MEASUREMENT_TACHO_MEASUREMENT(x) GetField(AXI_FAN_CONTROL_TACHO_MEASUREMENT,"TACHO_MEASUREMENT",x)
  `define DEFAULT_AXI_FAN_CONTROL_TACHO_MEASUREMENT_TACHO_MEASUREMENT GetResetValue(AXI_FAN_CONTROL_TACHO_MEASUREMENT,"TACHO_MEASUREMENT")
  `define UPDATE_AXI_FAN_CONTROL_TACHO_MEASUREMENT_TACHO_MEASUREMENT(x,y) UpdateField(AXI_FAN_CONTROL_TACHO_MEASUREMENT,"TACHO_MEASUREMENT",x,y)

  const reg_t AXI_FAN_CONTROL_TEMPERATURE = '{ 'h00c8, "TEMPERATURE" , '{
    "TEMPERATURE": '{ 31, 0, RO, 'h00000000 }}};
  `define SET_AXI_FAN_CONTROL_TEMPERATURE_TEMPERATURE(x) SetField(AXI_FAN_CONTROL_TEMPERATURE,"TEMPERATURE",x)
  `define GET_AXI_FAN_CONTROL_TEMPERATURE_TEMPERATURE(x) GetField(AXI_FAN_CONTROL_TEMPERATURE,"TEMPERATURE",x)
  `define DEFAULT_AXI_FAN_CONTROL_TEMPERATURE_TEMPERATURE GetResetValue(AXI_FAN_CONTROL_TEMPERATURE,"TEMPERATURE")
  `define UPDATE_AXI_FAN_CONTROL_TEMPERATURE_TEMPERATURE(x,y) UpdateField(AXI_FAN_CONTROL_TEMPERATURE,"TEMPERATURE",x,y)

  const reg_t AXI_FAN_CONTROL_TEMP_00_H = '{ 'h0100, "TEMP_00_H" , '{
    "TEMP_00_H": '{ 31, 0, RW, 0 }}};
  `define SET_AXI_FAN_CONTROL_TEMP_00_H_TEMP_00_H(x) SetField(AXI_FAN_CONTROL_TEMP_00_H,"TEMP_00_H",x)
  `define GET_AXI_FAN_CONTROL_TEMP_00_H_TEMP_00_H(x) GetField(AXI_FAN_CONTROL_TEMP_00_H,"TEMP_00_H",x)
  `define DEFAULT_AXI_FAN_CONTROL_TEMP_00_H_TEMP_00_H GetResetValue(AXI_FAN_CONTROL_TEMP_00_H,"TEMP_00_H")
  `define UPDATE_AXI_FAN_CONTROL_TEMP_00_H_TEMP_00_H(x,y) UpdateField(AXI_FAN_CONTROL_TEMP_00_H,"TEMP_00_H",x,y)

  const reg_t AXI_FAN_CONTROL_TEMP_25_L = '{ 'h0104, "TEMP_25_L" , '{
    "TEMP_25_L": '{ 31, 0, RW, 0 }}};
  `define SET_AXI_FAN_CONTROL_TEMP_25_L_TEMP_25_L(x) SetField(AXI_FAN_CONTROL_TEMP_25_L,"TEMP_25_L",x)
  `define GET_AXI_FAN_CONTROL_TEMP_25_L_TEMP_25_L(x) GetField(AXI_FAN_CONTROL_TEMP_25_L,"TEMP_25_L",x)
  `define DEFAULT_AXI_FAN_CONTROL_TEMP_25_L_TEMP_25_L GetResetValue(AXI_FAN_CONTROL_TEMP_25_L,"TEMP_25_L")
  `define UPDATE_AXI_FAN_CONTROL_TEMP_25_L_TEMP_25_L(x,y) UpdateField(AXI_FAN_CONTROL_TEMP_25_L,"TEMP_25_L",x,y)

  const reg_t AXI_FAN_CONTROL_TEMP_25_H = '{ 'h0108, "TEMP_25_H" , '{
    "TEMP_25_H": '{ 31, 0, RW, 0 }}};
  `define SET_AXI_FAN_CONTROL_TEMP_25_H_TEMP_25_H(x) SetField(AXI_FAN_CONTROL_TEMP_25_H,"TEMP_25_H",x)
  `define GET_AXI_FAN_CONTROL_TEMP_25_H_TEMP_25_H(x) GetField(AXI_FAN_CONTROL_TEMP_25_H,"TEMP_25_H",x)
  `define DEFAULT_AXI_FAN_CONTROL_TEMP_25_H_TEMP_25_H GetResetValue(AXI_FAN_CONTROL_TEMP_25_H,"TEMP_25_H")
  `define UPDATE_AXI_FAN_CONTROL_TEMP_25_H_TEMP_25_H(x,y) UpdateField(AXI_FAN_CONTROL_TEMP_25_H,"TEMP_25_H",x,y)

  const reg_t AXI_FAN_CONTROL_TEMP_50_L = '{ 'h010c, "TEMP_50_L" , '{
    "TEMP_50_L": '{ 31, 0, RW, 0 }}};
  `define SET_AXI_FAN_CONTROL_TEMP_50_L_TEMP_50_L(x) SetField(AXI_FAN_CONTROL_TEMP_50_L,"TEMP_50_L",x)
  `define GET_AXI_FAN_CONTROL_TEMP_50_L_TEMP_50_L(x) GetField(AXI_FAN_CONTROL_TEMP_50_L,"TEMP_50_L",x)
  `define DEFAULT_AXI_FAN_CONTROL_TEMP_50_L_TEMP_50_L GetResetValue(AXI_FAN_CONTROL_TEMP_50_L,"TEMP_50_L")
  `define UPDATE_AXI_FAN_CONTROL_TEMP_50_L_TEMP_50_L(x,y) UpdateField(AXI_FAN_CONTROL_TEMP_50_L,"TEMP_50_L",x,y)

  const reg_t AXI_FAN_CONTROL_TEMP_50_H = '{ 'h0110, "TEMP_50_H" , '{
    "TEMP_50_H": '{ 31, 0, RW, 0 }}};
  `define SET_AXI_FAN_CONTROL_TEMP_50_H_TEMP_50_H(x) SetField(AXI_FAN_CONTROL_TEMP_50_H,"TEMP_50_H",x)
  `define GET_AXI_FAN_CONTROL_TEMP_50_H_TEMP_50_H(x) GetField(AXI_FAN_CONTROL_TEMP_50_H,"TEMP_50_H",x)
  `define DEFAULT_AXI_FAN_CONTROL_TEMP_50_H_TEMP_50_H GetResetValue(AXI_FAN_CONTROL_TEMP_50_H,"TEMP_50_H")
  `define UPDATE_AXI_FAN_CONTROL_TEMP_50_H_TEMP_50_H(x,y) UpdateField(AXI_FAN_CONTROL_TEMP_50_H,"TEMP_50_H",x,y)

  const reg_t AXI_FAN_CONTROL_TEMP_75_L = '{ 'h0114, "TEMP_75_L" , '{
    "TEMP_75_L": '{ 31, 0, RW, 0 }}};
  `define SET_AXI_FAN_CONTROL_TEMP_75_L_TEMP_75_L(x) SetField(AXI_FAN_CONTROL_TEMP_75_L,"TEMP_75_L",x)
  `define GET_AXI_FAN_CONTROL_TEMP_75_L_TEMP_75_L(x) GetField(AXI_FAN_CONTROL_TEMP_75_L,"TEMP_75_L",x)
  `define DEFAULT_AXI_FAN_CONTROL_TEMP_75_L_TEMP_75_L GetResetValue(AXI_FAN_CONTROL_TEMP_75_L,"TEMP_75_L")
  `define UPDATE_AXI_FAN_CONTROL_TEMP_75_L_TEMP_75_L(x,y) UpdateField(AXI_FAN_CONTROL_TEMP_75_L,"TEMP_75_L",x,y)

  const reg_t AXI_FAN_CONTROL_TEMP_75_H = '{ 'h0118, "TEMP_75_H" , '{
    "TEMP_75_H": '{ 31, 0, RW, 0 }}};
  `define SET_AXI_FAN_CONTROL_TEMP_75_H_TEMP_75_H(x) SetField(AXI_FAN_CONTROL_TEMP_75_H,"TEMP_75_H",x)
  `define GET_AXI_FAN_CONTROL_TEMP_75_H_TEMP_75_H(x) GetField(AXI_FAN_CONTROL_TEMP_75_H,"TEMP_75_H",x)
  `define DEFAULT_AXI_FAN_CONTROL_TEMP_75_H_TEMP_75_H GetResetValue(AXI_FAN_CONTROL_TEMP_75_H,"TEMP_75_H")
  `define UPDATE_AXI_FAN_CONTROL_TEMP_75_H_TEMP_75_H(x,y) UpdateField(AXI_FAN_CONTROL_TEMP_75_H,"TEMP_75_H",x,y)

  const reg_t AXI_FAN_CONTROL_TEMP_100_L = '{ 'h011c, "TEMP_100_L" , '{
    "TEMP_100_L": '{ 31, 0, RW, 0 }}};
  `define SET_AXI_FAN_CONTROL_TEMP_100_L_TEMP_100_L(x) SetField(AXI_FAN_CONTROL_TEMP_100_L,"TEMP_100_L",x)
  `define GET_AXI_FAN_CONTROL_TEMP_100_L_TEMP_100_L(x) GetField(AXI_FAN_CONTROL_TEMP_100_L,"TEMP_100_L",x)
  `define DEFAULT_AXI_FAN_CONTROL_TEMP_100_L_TEMP_100_L GetResetValue(AXI_FAN_CONTROL_TEMP_100_L,"TEMP_100_L")
  `define UPDATE_AXI_FAN_CONTROL_TEMP_100_L_TEMP_100_L(x,y) UpdateField(AXI_FAN_CONTROL_TEMP_100_L,"TEMP_100_L",x,y)

  const reg_t AXI_FAN_CONTROL_TACHO_25 = '{ 'h0140, "TACHO_25" , '{
    "TACHO_25": '{ 31, 0, RW, 0 }}};
  `define SET_AXI_FAN_CONTROL_TACHO_25_TACHO_25(x) SetField(AXI_FAN_CONTROL_TACHO_25,"TACHO_25",x)
  `define GET_AXI_FAN_CONTROL_TACHO_25_TACHO_25(x) GetField(AXI_FAN_CONTROL_TACHO_25,"TACHO_25",x)
  `define DEFAULT_AXI_FAN_CONTROL_TACHO_25_TACHO_25 GetResetValue(AXI_FAN_CONTROL_TACHO_25,"TACHO_25")
  `define UPDATE_AXI_FAN_CONTROL_TACHO_25_TACHO_25(x,y) UpdateField(AXI_FAN_CONTROL_TACHO_25,"TACHO_25",x,y)

  const reg_t AXI_FAN_CONTROL_TACHO_50 = '{ 'h0144, "TACHO_50" , '{
    "TACHO_50": '{ 31, 0, RW, 0 }}};
  `define SET_AXI_FAN_CONTROL_TACHO_50_TACHO_50(x) SetField(AXI_FAN_CONTROL_TACHO_50,"TACHO_50",x)
  `define GET_AXI_FAN_CONTROL_TACHO_50_TACHO_50(x) GetField(AXI_FAN_CONTROL_TACHO_50,"TACHO_50",x)
  `define DEFAULT_AXI_FAN_CONTROL_TACHO_50_TACHO_50 GetResetValue(AXI_FAN_CONTROL_TACHO_50,"TACHO_50")
  `define UPDATE_AXI_FAN_CONTROL_TACHO_50_TACHO_50(x,y) UpdateField(AXI_FAN_CONTROL_TACHO_50,"TACHO_50",x,y)

  const reg_t AXI_FAN_CONTROL_TACHO_75 = '{ 'h0148, "TACHO_75" , '{
    "TACHO_75": '{ 31, 0, RW, 0 }}};
  `define SET_AXI_FAN_CONTROL_TACHO_75_TACHO_75(x) SetField(AXI_FAN_CONTROL_TACHO_75,"TACHO_75",x)
  `define GET_AXI_FAN_CONTROL_TACHO_75_TACHO_75(x) GetField(AXI_FAN_CONTROL_TACHO_75,"TACHO_75",x)
  `define DEFAULT_AXI_FAN_CONTROL_TACHO_75_TACHO_75 GetResetValue(AXI_FAN_CONTROL_TACHO_75,"TACHO_75")
  `define UPDATE_AXI_FAN_CONTROL_TACHO_75_TACHO_75(x,y) UpdateField(AXI_FAN_CONTROL_TACHO_75,"TACHO_75",x,y)

  const reg_t AXI_FAN_CONTROL_TACHO_100 = '{ 'h014c, "TACHO_100" , '{
    "TACHO_100": '{ 31, 0, RW, 0 }}};
  `define SET_AXI_FAN_CONTROL_TACHO_100_TACHO_100(x) SetField(AXI_FAN_CONTROL_TACHO_100,"TACHO_100",x)
  `define GET_AXI_FAN_CONTROL_TACHO_100_TACHO_100(x) GetField(AXI_FAN_CONTROL_TACHO_100,"TACHO_100",x)
  `define DEFAULT_AXI_FAN_CONTROL_TACHO_100_TACHO_100 GetResetValue(AXI_FAN_CONTROL_TACHO_100,"TACHO_100")
  `define UPDATE_AXI_FAN_CONTROL_TACHO_100_TACHO_100(x,y) UpdateField(AXI_FAN_CONTROL_TACHO_100,"TACHO_100",x,y)

  const reg_t AXI_FAN_CONTROL_TACHO_25_TOL = '{ 'h0150, "TACHO_25_TOL" , '{
    "TACHO_25_TOL": '{ 31, 0, RW, 0 }}};
  `define SET_AXI_FAN_CONTROL_TACHO_25_TOL_TACHO_25_TOL(x) SetField(AXI_FAN_CONTROL_TACHO_25_TOL,"TACHO_25_TOL",x)
  `define GET_AXI_FAN_CONTROL_TACHO_25_TOL_TACHO_25_TOL(x) GetField(AXI_FAN_CONTROL_TACHO_25_TOL,"TACHO_25_TOL",x)
  `define DEFAULT_AXI_FAN_CONTROL_TACHO_25_TOL_TACHO_25_TOL GetResetValue(AXI_FAN_CONTROL_TACHO_25_TOL,"TACHO_25_TOL")
  `define UPDATE_AXI_FAN_CONTROL_TACHO_25_TOL_TACHO_25_TOL(x,y) UpdateField(AXI_FAN_CONTROL_TACHO_25_TOL,"TACHO_25_TOL",x,y)

  const reg_t AXI_FAN_CONTROL_TACHO_50_TOL = '{ 'h0154, "TACHO_50_TOL" , '{
    "TACHO_50_TOL": '{ 31, 0, RW, 0 }}};
  `define SET_AXI_FAN_CONTROL_TACHO_50_TOL_TACHO_50_TOL(x) SetField(AXI_FAN_CONTROL_TACHO_50_TOL,"TACHO_50_TOL",x)
  `define GET_AXI_FAN_CONTROL_TACHO_50_TOL_TACHO_50_TOL(x) GetField(AXI_FAN_CONTROL_TACHO_50_TOL,"TACHO_50_TOL",x)
  `define DEFAULT_AXI_FAN_CONTROL_TACHO_50_TOL_TACHO_50_TOL GetResetValue(AXI_FAN_CONTROL_TACHO_50_TOL,"TACHO_50_TOL")
  `define UPDATE_AXI_FAN_CONTROL_TACHO_50_TOL_TACHO_50_TOL(x,y) UpdateField(AXI_FAN_CONTROL_TACHO_50_TOL,"TACHO_50_TOL",x,y)

  const reg_t AXI_FAN_CONTROL_TACHO_75_TOL = '{ 'h0158, "TACHO_75_TOL" , '{
    "TACHO_75_TOL": '{ 31, 0, RW, 0 }}};
  `define SET_AXI_FAN_CONTROL_TACHO_75_TOL_TACHO_75_TOL(x) SetField(AXI_FAN_CONTROL_TACHO_75_TOL,"TACHO_75_TOL",x)
  `define GET_AXI_FAN_CONTROL_TACHO_75_TOL_TACHO_75_TOL(x) GetField(AXI_FAN_CONTROL_TACHO_75_TOL,"TACHO_75_TOL",x)
  `define DEFAULT_AXI_FAN_CONTROL_TACHO_75_TOL_TACHO_75_TOL GetResetValue(AXI_FAN_CONTROL_TACHO_75_TOL,"TACHO_75_TOL")
  `define UPDATE_AXI_FAN_CONTROL_TACHO_75_TOL_TACHO_75_TOL(x,y) UpdateField(AXI_FAN_CONTROL_TACHO_75_TOL,"TACHO_75_TOL",x,y)

  const reg_t AXI_FAN_CONTROL_TACHO_100_TOL = '{ 'h015c, "TACHO_100_TOL" , '{
    "TACHO_100_TOL": '{ 31, 0, RW, 0 }}};
  `define SET_AXI_FAN_CONTROL_TACHO_100_TOL_TACHO_100_TOL(x) SetField(AXI_FAN_CONTROL_TACHO_100_TOL,"TACHO_100_TOL",x)
  `define GET_AXI_FAN_CONTROL_TACHO_100_TOL_TACHO_100_TOL(x) GetField(AXI_FAN_CONTROL_TACHO_100_TOL,"TACHO_100_TOL",x)
  `define DEFAULT_AXI_FAN_CONTROL_TACHO_100_TOL_TACHO_100_TOL GetResetValue(AXI_FAN_CONTROL_TACHO_100_TOL,"TACHO_100_TOL")
  `define UPDATE_AXI_FAN_CONTROL_TACHO_100_TOL_TACHO_100_TOL(x,y) UpdateField(AXI_FAN_CONTROL_TACHO_100_TOL,"TACHO_100_TOL",x,y)


endpackage
