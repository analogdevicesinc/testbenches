// ***************************************************************************
// ***************************************************************************
// Copyright 2024 (c) Analog Devices, Inc. All rights reserved.
//
// In this HDL repository, there are many different and unique modules, consisting
// of various HDL (Verilog or VHDL) components. The individual modules are
// developed independently, and may be accompanied by separate and unique license
// terms.
//
// The user should read each of these license terms, and understand the
// freedoms and responsabilities that he or she has by using this source/core.
//
// This core is distributed in the hope that it will be useful, but WITHOUT ANY
// WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR
// A PARTICULAR PURPOSE.
//
// Redistribution and use of source or resulting binaries, with or without modification
// of this file, are permitted under one of the following two license terms:
//
//   1. The GNU General Public License version 2 as published by the
//      Free Software Foundation, which can be found in the top level directory
//      of this repository (LICENSE_GPL2), and also online at:
//      <https://www.gnu.org/licenses/old-licenses/gpl-2.0.html>
//
// OR
//
//   2. An ADI specific BSD license, which can be found in the top level directory
//      of this repository (LICENSE_ADIBSD), and also on-line at:
//      https://github.com/analogdevicesinc/hdl/blob/master/LICENSE_ADIBSD
//      This will allow to generate bit files and not release the source code,
//      as long as it attaches to an ADI device.
//
// ***************************************************************************
// ***************************************************************************

`timescale 1ns/1ps

`include "utils.svh"

module system_tb();
  wire [3:0] quad_iso_adc_spi_cs;
  wire quad_iso_adc_spi_sclk;
  wire quad_iso_adc_spi_clk;
  wire [`NUM_OF_SDI-1:0] quad_iso_adc_spi_sdi;
  wire quad_iso_adc_spi_sdo;
  wire quad_iso_adc_irq;

  `TEST_PROGRAM test(
    .quad_iso_adc_irq(quad_iso_adc_irq),
    .quad_iso_adc_spi_sclk(quad_iso_adc_spi_sclk),
    .quad_iso_adc_spi_cs(quad_iso_adc_spi_cs),
    .quad_iso_adc_spi_clk(quad_iso_adc_spi_clk),
    .quad_iso_adc_spi_sdi(quad_iso_adc_spi_sdi));

  test_harness `TH (
    .quad_iso_adc_irq(quad_iso_adc_irq),
    .qadc_spi_cs(quad_iso_adc_spi_cs),
    .qadc_spi_sclk(quad_iso_adc_spi_sclk),
    .quad_iso_adc_spi_clk(quad_iso_adc_spi_clk),
    .qadc_spi_sdi(quad_iso_adc_spi_sdi),
    .qadc_spi_sdo(quad_iso_adc_spi_sdo));

endmodule
