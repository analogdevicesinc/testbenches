// ***************************************************************************
// ***************************************************************************
// Copyright (C) 2014 - 2025 Analog Devices, Inc. All rights reserved.
//
// In this HDL repository, there are many different and unique modules, consisting
// of various HDL (Verilog or VHDL) components. The individual modules are
// developed independently, and may be accompanied by separate and unique license
// terms.
//
// The user should read each of these license terms, and understand the
// freedoms and responsabilities that he or she has by using this source/core.
//
// This core is distributed in the hope that it will be useful, but WITHOUT ANY
// WARRANTY; without even the implied warranty of MERCHANTABILITY or FITNESS FOR
// A PARTICULAR PURPOSE.
//
// Redistribution and use of source or resulting binaries, with or without modification
// of this file, are permitted under one of the following two license terms:
//
//   1. The GNU General Public License version 2 as published by the
//      Free Software Foundation, which can be found in the top level directory
//      of this repository (LICENSE_GPL2), and also online at:
//      <https://www.gnu.org/licenses/old-licenses/gpl-2.0.html>
//
// OR
//
//   2. An ADI specific BSD license, which can be found in the top level directory
//      of this repository (LICENSE_ADIBSD), and also on-line at:
//      https://github.com/analogdevicesinc/hdl/blob/main/LICENSE_ADIBSD
//      This will allow to generate bit files and not release the source code,
//      as long as it attaches to an ADI device.
//
// ***************************************************************************
// ***************************************************************************
/* Auto generated Register Map */
/* Feb 07 14:25:05 2025 v0.4.1 */

`timescale 1ns/1ps

`ifndef _ADI_REGMAP_TDD_GEN_PKG_DEFINITIONS_SVH_
`define _ADI_REGMAP_TDD_GEN_PKG_DEFINITIONS_SVH_

// Help build VIP Interface parameters name
`define ADI_REGMAP_TDD_GEN_PKG_PARAM_IMPORT(n)  n``.inst.BURST_COUNT_WIDTH, \
  n``.inst.CHANNEL_COUNT, \
  n``.inst.DEFAULT_POLARITY, \
  n``.inst.ID, \
  n``.inst.REGISTER_WIDTH, \
  n``.inst.SYNC_COUNT_WIDTH, \
  n``.inst.SYNC_EXTERNAL, \
  n``.inst.SYNC_EXTERNAL_CDC, \
  n``.inst.SYNC_INTERNAL

`define ADI_REGMAP_TDD_GEN_PKG_PARAM_DECL int  BURST_COUNT_WIDTH, \
  CHANNEL_COUNT, \
  DEFAULT_POLARITY, \
  ID, \
  REGISTER_WIDTH, \
  SYNC_COUNT_WIDTH, \
  SYNC_EXTERNAL, \
  SYNC_EXTERNAL_CDC, \
  SYNC_INTERNAL

`define ADI_REGMAP_TDD_GEN_PKG_PARAM_ORDER  BURST_COUNT_WIDTH, \
  CHANNEL_COUNT, \
  DEFAULT_POLARITY, \
  ID, \
  REGISTER_WIDTH, \
  SYNC_COUNT_WIDTH, \
  SYNC_EXTERNAL, \
  SYNC_EXTERNAL_CDC, \
  SYNC_INTERNAL

`endif
